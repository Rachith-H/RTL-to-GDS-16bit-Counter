magic
tech sky130A
magscale 1 2
timestamp 1767199515
<< obsli1 >>
rect 1104 2159 11868 12529
<< obsm1 >>
rect 14 1436 12958 12560
<< metal2 >>
rect 1950 14346 2006 15146
rect 4526 14346 4582 15146
rect 7746 14346 7802 15146
rect 10322 14346 10378 15146
rect 12898 14346 12954 15146
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 8390 0 8446 800
rect 10966 0 11022 800
<< obsm2 >>
rect 20 14290 1894 14498
rect 2062 14290 4470 14498
rect 4638 14290 7690 14498
rect 7858 14290 10266 14498
rect 10434 14290 12842 14498
rect 20 856 12952 14290
rect 130 711 2538 856
rect 2706 711 5114 856
rect 5282 711 8334 856
rect 8502 711 10910 856
rect 11078 711 12952 856
<< metal3 >>
rect 0 14288 800 14408
rect 12202 12248 13002 12368
rect 0 11568 800 11688
rect 12202 9528 13002 9648
rect 0 8848 800 8968
rect 12202 6128 13002 6248
rect 0 5448 800 5568
rect 12202 3408 13002 3528
rect 0 2728 800 2848
rect 12202 688 13002 808
<< obsm3 >>
rect 880 14208 12202 14378
rect 800 12448 12202 14208
rect 800 12168 12122 12448
rect 800 11768 12202 12168
rect 880 11488 12202 11768
rect 800 9728 12202 11488
rect 800 9448 12122 9728
rect 800 9048 12202 9448
rect 880 8768 12202 9048
rect 800 6328 12202 8768
rect 800 6048 12122 6328
rect 800 5648 12202 6048
rect 880 5368 12202 5648
rect 800 3608 12202 5368
rect 800 3328 12122 3608
rect 800 2928 12202 3328
rect 880 2648 12202 2928
rect 800 888 12202 2648
rect 800 715 12122 888
<< metal4 >>
rect 2289 2128 2609 12560
rect 2949 2128 3269 12560
rect 4980 2128 5300 12560
rect 5640 2128 5960 12560
rect 7671 2128 7991 12560
rect 8331 2128 8651 12560
rect 10362 2128 10682 12560
rect 11022 2128 11342 12560
<< obsm4 >>
rect 6867 3435 7591 7037
rect 8071 3435 8251 7037
rect 8731 3435 9693 7037
<< metal5 >>
rect 1056 11720 11916 12040
rect 1056 11060 11916 11380
rect 1056 9136 11916 9456
rect 1056 8476 11916 8796
rect 1056 6552 11916 6872
rect 1056 5892 11916 6212
rect 1056 3968 11916 4288
rect 1056 3308 11916 3628
<< labels >>
rlabel metal4 s 2949 2128 3269 12560 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 5640 2128 5960 12560 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8331 2128 8651 12560 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11022 2128 11342 12560 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3968 11916 4288 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6552 11916 6872 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9136 11916 9456 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 11720 11916 12040 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2289 2128 2609 12560 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4980 2128 5300 12560 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7671 2128 7991 12560 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 10362 2128 10682 12560 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3308 11916 3628 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5892 11916 6212 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8476 11916 8796 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11060 11916 11380 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 12202 3408 13002 3528 6 clk
port 3 nsew signal input
rlabel metal2 s 12898 14346 12954 15146 6 count[0]
port 4 nsew signal output
rlabel metal2 s 7746 14346 7802 15146 6 count[10]
port 5 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 count[11]
port 6 nsew signal output
rlabel metal3 s 12202 12248 13002 12368 6 count[12]
port 7 nsew signal output
rlabel metal3 s 12202 688 13002 808 6 count[13]
port 8 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 count[14]
port 9 nsew signal output
rlabel metal2 s 4526 14346 4582 15146 6 count[15]
port 10 nsew signal output
rlabel metal2 s 18 0 74 800 6 count[1]
port 11 nsew signal output
rlabel metal2 s 1950 14346 2006 15146 6 count[2]
port 12 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 count[3]
port 13 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 count[4]
port 14 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 count[5]
port 15 nsew signal output
rlabel metal3 s 12202 9528 13002 9648 6 count[6]
port 16 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 count[7]
port 17 nsew signal output
rlabel metal2 s 10322 14346 10378 15146 6 count[8]
port 18 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 count[9]
port 19 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 ctrl
port 20 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 en
port 21 nsew signal input
rlabel metal3 s 12202 6128 13002 6248 6 rst
port 22 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 13002 15146
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 707786
string GDS_FILE /openlane/designs/counter_up_dwn/runs/RUN_2025.12.31_16.42.11/results/signoff/counter_up_dwn.magic.gds
string GDS_START 289490
<< end >>

