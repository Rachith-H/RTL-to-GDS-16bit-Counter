VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter_up_dwn
  CLASS BLOCK ;
  FOREIGN counter_up_dwn ;
  ORIGIN 0.000 0.000 ;
  SIZE 65.010 BY 75.730 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.745 10.640 16.345 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.200 10.640 29.800 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.655 10.640 43.255 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.110 10.640 56.710 62.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.840 59.580 21.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 32.760 59.580 34.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 45.680 59.580 47.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 58.600 59.580 60.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.445 10.640 13.045 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.900 10.640 26.500 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.355 10.640 39.955 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.810 10.640 53.410 62.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 16.540 59.580 18.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 29.460 59.580 31.060 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 42.380 59.580 43.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 55.300 59.580 56.900 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 61.010 17.040 65.010 17.640 ;
    END
  END clk
  PIN count[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 71.730 64.770 75.730 ;
    END
  END count[0]
  PIN count[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.730 71.730 39.010 75.730 ;
    END
  END count[10]
  PIN count[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END count[11]
  PIN count[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 61.010 61.240 65.010 61.840 ;
    END
  END count[12]
  PIN count[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 61.010 3.440 65.010 4.040 ;
    END
  END count[13]
  PIN count[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END count[14]
  PIN count[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 71.730 22.910 75.730 ;
    END
  END count[15]
  PIN count[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END count[1]
  PIN count[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 9.750 71.730 10.030 75.730 ;
    END
  END count[2]
  PIN count[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END count[3]
  PIN count[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END count[4]
  PIN count[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END count[5]
  PIN count[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 61.010 47.640 65.010 48.240 ;
    END
  END count[6]
  PIN count[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END count[7]
  PIN count[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 51.610 71.730 51.890 75.730 ;
    END
  END count[8]
  PIN count[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END count[9]
  PIN ctrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END ctrl
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END en
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 61.010 30.640 65.010 31.240 ;
    END
  END rst
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 59.340 62.645 ;
      LAYER met1 ;
        RECT 0.070 7.180 64.790 62.800 ;
      LAYER met2 ;
        RECT 0.100 71.450 9.470 72.490 ;
        RECT 10.310 71.450 22.350 72.490 ;
        RECT 23.190 71.450 38.450 72.490 ;
        RECT 39.290 71.450 51.330 72.490 ;
        RECT 52.170 71.450 64.210 72.490 ;
        RECT 0.100 4.280 64.760 71.450 ;
        RECT 0.650 3.555 12.690 4.280 ;
        RECT 13.530 3.555 25.570 4.280 ;
        RECT 26.410 3.555 41.670 4.280 ;
        RECT 42.510 3.555 54.550 4.280 ;
        RECT 55.390 3.555 64.760 4.280 ;
      LAYER met3 ;
        RECT 4.400 71.040 61.010 71.890 ;
        RECT 4.000 62.240 61.010 71.040 ;
        RECT 4.000 60.840 60.610 62.240 ;
        RECT 4.000 58.840 61.010 60.840 ;
        RECT 4.400 57.440 61.010 58.840 ;
        RECT 4.000 48.640 61.010 57.440 ;
        RECT 4.000 47.240 60.610 48.640 ;
        RECT 4.000 45.240 61.010 47.240 ;
        RECT 4.400 43.840 61.010 45.240 ;
        RECT 4.000 31.640 61.010 43.840 ;
        RECT 4.000 30.240 60.610 31.640 ;
        RECT 4.000 28.240 61.010 30.240 ;
        RECT 4.400 26.840 61.010 28.240 ;
        RECT 4.000 18.040 61.010 26.840 ;
        RECT 4.000 16.640 60.610 18.040 ;
        RECT 4.000 14.640 61.010 16.640 ;
        RECT 4.400 13.240 61.010 14.640 ;
        RECT 4.000 4.440 61.010 13.240 ;
        RECT 4.000 3.575 60.610 4.440 ;
      LAYER met4 ;
        RECT 34.335 17.175 37.955 35.185 ;
        RECT 40.355 17.175 41.255 35.185 ;
        RECT 43.655 17.175 48.465 35.185 ;
  END
END counter_up_dwn
END LIBRARY

