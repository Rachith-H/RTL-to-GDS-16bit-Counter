magic
tech sky130A
magscale 1 2
timestamp 1767199513
<< viali >>
rect 2973 12393 3007 12427
rect 4721 12393 4755 12427
rect 10609 12393 10643 12427
rect 11253 12393 11287 12427
rect 8033 12325 8067 12359
rect 10149 12257 10183 12291
rect 1409 12189 1443 12223
rect 2145 12189 2179 12223
rect 11069 12189 11103 12223
rect 3249 12121 3283 12155
rect 4997 12121 5031 12155
rect 8217 12121 8251 12155
rect 10517 12121 10551 12155
rect 1593 12053 1627 12087
rect 2789 12053 2823 12087
rect 9597 12053 9631 12087
rect 10609 11849 10643 11883
rect 11253 11849 11287 11883
rect 1777 11781 1811 11815
rect 9137 11781 9171 11815
rect 10977 11781 11011 11815
rect 1409 11713 1443 11747
rect 2421 11713 2455 11747
rect 2789 11713 2823 11747
rect 5089 11713 5123 11747
rect 5733 11713 5767 11747
rect 6745 11713 6779 11747
rect 8401 11713 8435 11747
rect 2329 11645 2363 11679
rect 2697 11645 2731 11679
rect 3065 11645 3099 11679
rect 4537 11645 4571 11679
rect 4813 11645 4847 11679
rect 4997 11645 5031 11679
rect 8493 11645 8527 11679
rect 8769 11645 8803 11679
rect 8861 11645 8895 11679
rect 2145 11509 2179 11543
rect 5457 11509 5491 11543
rect 5549 11509 5583 11543
rect 6653 11509 6687 11543
rect 3249 11305 3283 11339
rect 4629 11305 4663 11339
rect 5168 11305 5202 11339
rect 8493 11305 8527 11339
rect 9781 11305 9815 11339
rect 2881 11169 2915 11203
rect 3157 11169 3191 11203
rect 4905 11169 4939 11203
rect 6745 11169 6779 11203
rect 9505 11169 9539 11203
rect 3525 11101 3559 11135
rect 4353 11101 4387 11135
rect 4721 11101 4755 11135
rect 8769 11101 8803 11135
rect 9689 11101 9723 11135
rect 10149 11101 10183 11135
rect 3249 11033 3283 11067
rect 7021 11033 7055 11067
rect 8677 11033 8711 11067
rect 1409 10965 1443 10999
rect 3433 10965 3467 10999
rect 3801 10965 3835 10999
rect 6653 10965 6687 10999
rect 8953 10965 8987 10999
rect 9965 10965 9999 10999
rect 2421 10761 2455 10795
rect 3985 10761 4019 10795
rect 5457 10761 5491 10795
rect 5825 10761 5859 10795
rect 6561 10761 6595 10795
rect 6929 10761 6963 10795
rect 7113 10761 7147 10795
rect 8493 10761 8527 10795
rect 11345 10761 11379 10795
rect 7665 10693 7699 10727
rect 7757 10693 7791 10727
rect 9873 10693 9907 10727
rect 2513 10625 2547 10659
rect 2761 10625 2795 10659
rect 3341 10625 3375 10659
rect 3433 10625 3467 10659
rect 3617 10625 3651 10659
rect 3709 10625 3743 10659
rect 3801 10625 3835 10659
rect 4353 10625 4387 10659
rect 4537 10625 4571 10659
rect 4813 10625 4847 10659
rect 6469 10625 6503 10659
rect 6653 10625 6687 10659
rect 6745 10625 6779 10659
rect 7021 10625 7055 10659
rect 7389 10625 7423 10659
rect 8033 10625 8067 10659
rect 8217 10625 8251 10659
rect 8309 10625 8343 10659
rect 8401 10625 8435 10659
rect 8585 10625 8619 10659
rect 2927 10557 2961 10591
rect 4261 10557 4295 10591
rect 4445 10557 4479 10591
rect 5917 10557 5951 10591
rect 6101 10557 6135 10591
rect 7297 10557 7331 10591
rect 9597 10557 9631 10591
rect 3065 10489 3099 10523
rect 4077 10489 4111 10523
rect 5089 10489 5123 10523
rect 7849 10489 7883 10523
rect 6745 10421 6779 10455
rect 2789 10217 2823 10251
rect 2973 10217 3007 10251
rect 3433 10217 3467 10251
rect 4169 10217 4203 10251
rect 4997 10217 5031 10251
rect 5917 10217 5951 10251
rect 7205 10217 7239 10251
rect 7665 10217 7699 10251
rect 10241 10217 10275 10251
rect 10885 10217 10919 10251
rect 3801 10149 3835 10183
rect 4261 10081 4295 10115
rect 5549 10081 5583 10115
rect 9689 10081 9723 10115
rect 2421 10013 2455 10047
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 3341 10013 3375 10047
rect 3525 10013 3559 10047
rect 3985 10013 4019 10047
rect 4905 10013 4939 10047
rect 5641 10013 5675 10047
rect 7389 10013 7423 10047
rect 7573 10013 7607 10047
rect 7665 10013 7699 10047
rect 7849 10013 7883 10047
rect 10977 10013 11011 10047
rect 2605 9945 2639 9979
rect 9873 9945 9907 9979
rect 11161 9945 11195 9979
rect 9781 9877 9815 9911
rect 11437 9877 11471 9911
rect 2421 9605 2455 9639
rect 9321 9605 9355 9639
rect 9505 9605 9539 9639
rect 2605 9537 2639 9571
rect 8861 9537 8895 9571
rect 9781 9537 9815 9571
rect 9965 9537 9999 9571
rect 8953 9469 8987 9503
rect 9229 9469 9263 9503
rect 2789 9333 2823 9367
rect 9689 9333 9723 9367
rect 9873 9333 9907 9367
rect 3249 9129 3283 9163
rect 6653 9129 6687 9163
rect 10057 9129 10091 9163
rect 8677 9061 8711 9095
rect 4905 8993 4939 9027
rect 8769 8993 8803 9027
rect 9689 8993 9723 9027
rect 9873 8993 9907 9027
rect 10333 8993 10367 9027
rect 1409 8925 1443 8959
rect 3065 8925 3099 8959
rect 3341 8925 3375 8959
rect 3433 8925 3467 8959
rect 3617 8925 3651 8959
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 4261 8925 4295 8959
rect 6929 8925 6963 8959
rect 8493 8925 8527 8959
rect 8953 8925 8987 8959
rect 9321 8925 9355 8959
rect 9413 8925 9447 8959
rect 10148 8903 10182 8937
rect 10241 8925 10275 8959
rect 10425 8925 10459 8959
rect 2053 8857 2087 8891
rect 2421 8857 2455 8891
rect 4537 8857 4571 8891
rect 4629 8857 4663 8891
rect 5181 8857 5215 8891
rect 9781 8857 9815 8891
rect 9873 8857 9907 8891
rect 1593 8789 1627 8823
rect 2881 8789 2915 8823
rect 3617 8789 3651 8823
rect 7021 8789 7055 8823
rect 8309 8789 8343 8823
rect 3157 8585 3191 8619
rect 3801 8585 3835 8619
rect 4721 8585 4755 8619
rect 5181 8585 5215 8619
rect 6009 8585 6043 8619
rect 11345 8585 11379 8619
rect 6653 8517 6687 8551
rect 8677 8517 8711 8551
rect 2053 8449 2087 8483
rect 2789 8449 2823 8483
rect 3065 8449 3099 8483
rect 3249 8449 3283 8483
rect 3525 8449 3559 8483
rect 3617 8449 3651 8483
rect 5365 8449 5399 8483
rect 5917 8449 5951 8483
rect 6377 8449 6411 8483
rect 8769 8449 8803 8483
rect 9045 8449 9079 8483
rect 9597 8449 9631 8483
rect 2145 8381 2179 8415
rect 3801 8381 3835 8415
rect 4445 8381 4479 8415
rect 4629 8381 4663 8415
rect 8953 8381 8987 8415
rect 9873 8381 9907 8415
rect 2421 8313 2455 8347
rect 2881 8313 2915 8347
rect 5089 8313 5123 8347
rect 8125 8313 8159 8347
rect 9413 8313 9447 8347
rect 5733 8041 5767 8075
rect 8953 8041 8987 8075
rect 10425 8041 10459 8075
rect 10885 8041 10919 8075
rect 10333 7973 10367 8007
rect 2329 7905 2363 7939
rect 8125 7905 8159 7939
rect 9229 7905 9263 7939
rect 9689 7905 9723 7939
rect 9873 7905 9907 7939
rect 3433 7837 3467 7871
rect 3617 7837 3651 7871
rect 8309 7837 8343 7871
rect 8585 7837 8619 7871
rect 9321 7837 9355 7871
rect 10609 7837 10643 7871
rect 10977 7837 11011 7871
rect 1777 7769 1811 7803
rect 7021 7769 7055 7803
rect 3525 7701 3559 7735
rect 7573 7701 7607 7735
rect 9965 7701 9999 7735
rect 3065 7497 3099 7531
rect 4261 7429 4295 7463
rect 3249 7361 3283 7395
rect 3709 7361 3743 7395
rect 8125 7361 8159 7395
rect 3433 7293 3467 7327
rect 3801 7293 3835 7327
rect 4077 7293 4111 7327
rect 4537 7157 4571 7191
rect 6837 7157 6871 7191
rect 3617 6953 3651 6987
rect 7113 6953 7147 6987
rect 7297 6953 7331 6987
rect 7665 6953 7699 6987
rect 1869 6817 1903 6851
rect 2145 6817 2179 6851
rect 6561 6817 6595 6851
rect 9965 6817 9999 6851
rect 10057 6817 10091 6851
rect 1777 6749 1811 6783
rect 3065 6749 3099 6783
rect 3341 6749 3375 6783
rect 3433 6749 3467 6783
rect 3617 6749 3651 6783
rect 5825 6749 5859 6783
rect 6101 6749 6135 6783
rect 6653 6749 6687 6783
rect 6929 6749 6963 6783
rect 7021 6749 7055 6783
rect 7573 6749 7607 6783
rect 7757 6749 7791 6783
rect 8493 6749 8527 6783
rect 8677 6749 8711 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 9413 6749 9447 6783
rect 9873 6749 9907 6783
rect 10149 6749 10183 6783
rect 3249 6681 3283 6715
rect 5917 6681 5951 6715
rect 7481 6681 7515 6715
rect 3163 6613 3197 6647
rect 6285 6613 6319 6647
rect 6377 6613 6411 6647
rect 7281 6613 7315 6647
rect 8585 6613 8619 6647
rect 9597 6613 9631 6647
rect 9689 6613 9723 6647
rect 3341 6409 3375 6443
rect 3893 6409 3927 6443
rect 5181 6409 5215 6443
rect 5825 6409 5859 6443
rect 7113 6409 7147 6443
rect 7573 6409 7607 6443
rect 8309 6409 8343 6443
rect 9413 6409 9447 6443
rect 4905 6341 4939 6375
rect 6745 6341 6779 6375
rect 9781 6341 9815 6375
rect 2145 6273 2179 6307
rect 4169 6273 4203 6307
rect 4353 6273 4387 6307
rect 4530 6273 4564 6307
rect 4629 6273 4663 6307
rect 4813 6273 4847 6307
rect 5089 6273 5123 6307
rect 5181 6273 5215 6307
rect 5273 6273 5307 6307
rect 5825 6273 5859 6307
rect 6469 6273 6503 6307
rect 6653 6273 6687 6307
rect 6929 6273 6963 6307
rect 7205 6273 7239 6307
rect 7389 6273 7423 6307
rect 7489 6271 7523 6305
rect 7665 6273 7699 6307
rect 7941 6273 7975 6307
rect 8125 6273 8159 6307
rect 8585 6273 8619 6307
rect 9229 6273 9263 6307
rect 2237 6205 2271 6239
rect 3893 6205 3927 6239
rect 7297 6205 7331 6239
rect 7849 6205 7883 6239
rect 8677 6205 8711 6239
rect 9045 6205 9079 6239
rect 9505 6205 9539 6239
rect 2513 6137 2547 6171
rect 2973 6137 3007 6171
rect 4077 6137 4111 6171
rect 5438 6137 5472 6171
rect 3341 6069 3375 6103
rect 3525 6069 3559 6103
rect 4445 6069 4479 6103
rect 4813 6069 4847 6103
rect 5549 6069 5583 6103
rect 5641 6069 5675 6103
rect 6561 6069 6595 6103
rect 8953 6069 8987 6103
rect 11253 6069 11287 6103
rect 4445 5865 4479 5899
rect 8217 5865 8251 5899
rect 8953 5865 8987 5899
rect 9321 5865 9355 5899
rect 10885 5865 10919 5899
rect 8769 5797 8803 5831
rect 11161 5797 11195 5831
rect 1961 5729 1995 5763
rect 4169 5729 4203 5763
rect 5273 5729 5307 5763
rect 5457 5729 5491 5763
rect 9045 5729 9079 5763
rect 9413 5729 9447 5763
rect 9781 5729 9815 5763
rect 2237 5661 2271 5695
rect 4077 5661 4111 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 5089 5661 5123 5695
rect 5549 5661 5583 5695
rect 8033 5661 8067 5695
rect 8309 5661 8343 5695
rect 8401 5661 8435 5695
rect 8493 5661 8527 5695
rect 8953 5661 8987 5695
rect 9873 5661 9907 5695
rect 10977 5661 11011 5695
rect 11437 5661 11471 5695
rect 5181 5593 5215 5627
rect 2881 5525 2915 5559
rect 4537 5525 4571 5559
rect 5273 5525 5307 5559
rect 10057 5525 10091 5559
rect 2421 5321 2455 5355
rect 4721 5321 4755 5355
rect 6561 5321 6595 5355
rect 8769 5321 8803 5355
rect 1409 5253 1443 5287
rect 1777 5253 1811 5287
rect 2329 5253 2363 5287
rect 4537 5185 4571 5219
rect 4721 5185 4755 5219
rect 6469 5185 6503 5219
rect 8953 5185 8987 5219
rect 9321 5185 9355 5219
rect 9413 5185 9447 5219
rect 9505 5185 9539 5219
rect 2513 5117 2547 5151
rect 9689 5117 9723 5151
rect 9597 5049 9631 5083
rect 1961 4981 1995 5015
rect 9229 4981 9263 5015
rect 5641 4777 5675 4811
rect 9413 4777 9447 4811
rect 7481 4709 7515 4743
rect 4445 4641 4479 4675
rect 7021 4641 7055 4675
rect 7849 4641 7883 4675
rect 9045 4641 9079 4675
rect 10057 4641 10091 4675
rect 2145 4573 2179 4607
rect 4905 4573 4939 4607
rect 6285 4573 6319 4607
rect 7113 4573 7147 4607
rect 7941 4573 7975 4607
rect 9137 4573 9171 4607
rect 9965 4573 9999 4607
rect 4813 4505 4847 4539
rect 1961 4437 1995 4471
rect 4721 4437 4755 4471
rect 7573 4437 7607 4471
rect 9597 4437 9631 4471
rect 4537 4233 4571 4267
rect 1869 4165 1903 4199
rect 1593 4097 1627 4131
rect 3709 4097 3743 4131
rect 4997 4097 5031 4131
rect 5457 4097 5491 4131
rect 5733 4097 5767 4131
rect 8769 4097 8803 4131
rect 3801 4029 3835 4063
rect 4261 4029 4295 4063
rect 4445 4029 4479 4063
rect 4077 3961 4111 3995
rect 4905 3961 4939 3995
rect 3341 3893 3375 3927
rect 5181 3893 5215 3927
rect 5365 3893 5399 3927
rect 5641 3893 5675 3927
rect 8861 3893 8895 3927
rect 3525 3689 3559 3723
rect 4905 3621 4939 3655
rect 8953 3621 8987 3655
rect 2053 3553 2087 3587
rect 6285 3553 6319 3587
rect 9505 3553 9539 3587
rect 1777 3485 1811 3519
rect 2237 3485 2271 3519
rect 2973 3485 3007 3519
rect 3617 3485 3651 3519
rect 6193 3485 6227 3519
rect 8585 3485 8619 3519
rect 9321 3485 9355 3519
rect 9413 3485 9447 3519
rect 1409 3417 1443 3451
rect 6561 3417 6595 3451
rect 2329 3349 2363 3383
rect 2697 3349 2731 3383
rect 2789 3349 2823 3383
rect 8033 3349 8067 3383
rect 8401 3349 8435 3383
rect 6653 3145 6687 3179
rect 7389 3145 7423 3179
rect 9505 3145 9539 3179
rect 3893 3077 3927 3111
rect 4445 3077 4479 3111
rect 7297 3077 7331 3111
rect 1685 3009 1719 3043
rect 3985 3009 4019 3043
rect 4169 3009 4203 3043
rect 6837 3009 6871 3043
rect 7764 3009 7798 3043
rect 10977 3009 11011 3043
rect 1961 2941 1995 2975
rect 3709 2941 3743 2975
rect 6193 2941 6227 2975
rect 7573 2941 7607 2975
rect 8033 2941 8067 2975
rect 6929 2873 6963 2907
rect 11069 2805 11103 2839
rect 7389 2601 7423 2635
rect 3985 2465 4019 2499
rect 5733 2465 5767 2499
rect 6009 2465 6043 2499
rect 1777 2397 1811 2431
rect 2881 2397 2915 2431
rect 7297 2397 7331 2431
rect 9045 2397 9079 2431
rect 10977 2397 11011 2431
rect 1409 2329 1443 2363
rect 6377 2329 6411 2363
rect 6745 2329 6779 2363
rect 2605 2261 2639 2295
rect 9137 2261 9171 2295
rect 11069 2261 11103 2295
<< metal1 >>
rect 1104 12538 11868 12560
rect 1104 12486 2295 12538
rect 2347 12486 2359 12538
rect 2411 12486 2423 12538
rect 2475 12486 2487 12538
rect 2539 12486 2551 12538
rect 2603 12486 4986 12538
rect 5038 12486 5050 12538
rect 5102 12486 5114 12538
rect 5166 12486 5178 12538
rect 5230 12486 5242 12538
rect 5294 12486 7677 12538
rect 7729 12486 7741 12538
rect 7793 12486 7805 12538
rect 7857 12486 7869 12538
rect 7921 12486 7933 12538
rect 7985 12486 10368 12538
rect 10420 12486 10432 12538
rect 10484 12486 10496 12538
rect 10548 12486 10560 12538
rect 10612 12486 10624 12538
rect 10676 12486 11868 12538
rect 1104 12464 11868 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 2961 12427 3019 12433
rect 2961 12424 2973 12427
rect 2004 12396 2973 12424
rect 2004 12384 2010 12396
rect 2961 12393 2973 12396
rect 3007 12393 3019 12427
rect 2961 12387 3019 12393
rect 4706 12384 4712 12436
rect 4764 12384 4770 12436
rect 10226 12384 10232 12436
rect 10284 12424 10290 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 10284 12396 10609 12424
rect 10284 12384 10290 12396
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 10597 12387 10655 12393
rect 11238 12384 11244 12436
rect 11296 12384 11302 12436
rect 8018 12316 8024 12368
rect 8076 12316 8082 12368
rect 2222 12248 2228 12300
rect 2280 12288 2286 12300
rect 2280 12260 2774 12288
rect 2280 12248 2286 12260
rect 1394 12180 1400 12232
rect 1452 12180 1458 12232
rect 1854 12180 1860 12232
rect 1912 12220 1918 12232
rect 2133 12223 2191 12229
rect 2133 12220 2145 12223
rect 1912 12192 2145 12220
rect 1912 12180 1918 12192
rect 2133 12189 2145 12192
rect 2179 12189 2191 12223
rect 2746 12220 2774 12260
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 10134 12288 10140 12300
rect 4764 12260 10140 12288
rect 4764 12248 4770 12260
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 8662 12220 8668 12232
rect 2746 12192 8668 12220
rect 2133 12183 2191 12189
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12220 11115 12223
rect 11422 12220 11428 12232
rect 11103 12192 11428 12220
rect 11103 12189 11115 12192
rect 11057 12183 11115 12189
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 3237 12155 3295 12161
rect 3237 12121 3249 12155
rect 3283 12152 3295 12155
rect 3418 12152 3424 12164
rect 3283 12124 3424 12152
rect 3283 12121 3295 12124
rect 3237 12115 3295 12121
rect 3418 12112 3424 12124
rect 3476 12112 3482 12164
rect 4982 12112 4988 12164
rect 5040 12112 5046 12164
rect 8110 12112 8116 12164
rect 8168 12152 8174 12164
rect 8205 12155 8263 12161
rect 8205 12152 8217 12155
rect 8168 12124 8217 12152
rect 8168 12112 8174 12124
rect 8205 12121 8217 12124
rect 8251 12121 8263 12155
rect 10505 12155 10563 12161
rect 10505 12152 10517 12155
rect 8205 12115 8263 12121
rect 8312 12124 10517 12152
rect 1578 12044 1584 12096
rect 1636 12044 1642 12096
rect 2774 12044 2780 12096
rect 2832 12044 2838 12096
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8312 12084 8340 12124
rect 10505 12121 10517 12124
rect 10551 12121 10563 12155
rect 10505 12115 10563 12121
rect 8076 12056 8340 12084
rect 8076 12044 8082 12056
rect 9030 12044 9036 12096
rect 9088 12084 9094 12096
rect 9585 12087 9643 12093
rect 9585 12084 9597 12087
rect 9088 12056 9597 12084
rect 9088 12044 9094 12056
rect 9585 12053 9597 12056
rect 9631 12053 9643 12087
rect 9585 12047 9643 12053
rect 1104 11994 11868 12016
rect 1104 11942 2955 11994
rect 3007 11942 3019 11994
rect 3071 11942 3083 11994
rect 3135 11942 3147 11994
rect 3199 11942 3211 11994
rect 3263 11942 5646 11994
rect 5698 11942 5710 11994
rect 5762 11942 5774 11994
rect 5826 11942 5838 11994
rect 5890 11942 5902 11994
rect 5954 11942 8337 11994
rect 8389 11942 8401 11994
rect 8453 11942 8465 11994
rect 8517 11942 8529 11994
rect 8581 11942 8593 11994
rect 8645 11942 11028 11994
rect 11080 11942 11092 11994
rect 11144 11942 11156 11994
rect 11208 11942 11220 11994
rect 11272 11942 11284 11994
rect 11336 11942 11868 11994
rect 1104 11920 11868 11942
rect 2222 11840 2228 11892
rect 2280 11840 2286 11892
rect 2774 11840 2780 11892
rect 2832 11840 2838 11892
rect 3694 11880 3700 11892
rect 2976 11852 3700 11880
rect 1765 11815 1823 11821
rect 1765 11781 1777 11815
rect 1811 11812 1823 11815
rect 2240 11812 2268 11840
rect 1811 11784 2268 11812
rect 1811 11781 1823 11784
rect 1765 11775 1823 11781
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 2792 11753 2820 11840
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11713 2467 11747
rect 2409 11707 2467 11713
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11645 2375 11679
rect 2317 11639 2375 11645
rect 2130 11500 2136 11552
rect 2188 11500 2194 11552
rect 2332 11540 2360 11639
rect 2424 11608 2452 11707
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 2976 11676 3004 11852
rect 3694 11840 3700 11852
rect 3752 11840 3758 11892
rect 4982 11840 4988 11892
rect 5040 11840 5046 11892
rect 9030 11880 9036 11892
rect 8680 11852 9036 11880
rect 4062 11772 4068 11824
rect 4120 11772 4126 11824
rect 5000 11812 5028 11840
rect 5994 11812 6000 11824
rect 5000 11784 6000 11812
rect 5000 11744 5028 11784
rect 5994 11772 6000 11784
rect 6052 11772 6058 11824
rect 5077 11747 5135 11753
rect 5077 11744 5089 11747
rect 5000 11716 5089 11744
rect 5077 11713 5089 11716
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 5721 11747 5779 11753
rect 5721 11744 5733 11747
rect 5408 11716 5733 11744
rect 5408 11704 5414 11716
rect 5721 11713 5733 11716
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 8294 11744 8300 11756
rect 6779 11716 8300 11744
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 8294 11704 8300 11716
rect 8352 11704 8358 11756
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11713 8447 11747
rect 8389 11707 8447 11713
rect 2731 11648 3004 11676
rect 3053 11679 3111 11685
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 3053 11645 3065 11679
rect 3099 11676 3111 11679
rect 3099 11648 3464 11676
rect 3099 11645 3111 11648
rect 3053 11639 3111 11645
rect 2424 11580 3280 11608
rect 3252 11552 3280 11580
rect 3436 11552 3464 11648
rect 4522 11636 4528 11688
rect 4580 11636 4586 11688
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11645 4859 11679
rect 4801 11639 4859 11645
rect 4816 11608 4844 11639
rect 4890 11636 4896 11688
rect 4948 11676 4954 11688
rect 4985 11679 5043 11685
rect 4985 11676 4997 11679
rect 4948 11648 4997 11676
rect 4948 11636 4954 11648
rect 4985 11645 4997 11648
rect 5031 11645 5043 11679
rect 4985 11639 5043 11645
rect 5534 11636 5540 11688
rect 5592 11636 5598 11688
rect 5552 11608 5580 11636
rect 4816 11580 5580 11608
rect 8404 11608 8432 11707
rect 8481 11679 8539 11685
rect 8481 11645 8493 11679
rect 8527 11676 8539 11679
rect 8680 11676 8708 11852
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10597 11883 10655 11889
rect 10597 11880 10609 11883
rect 10192 11852 10609 11880
rect 10192 11840 10198 11852
rect 10597 11849 10609 11852
rect 10643 11880 10655 11883
rect 11241 11883 11299 11889
rect 10643 11852 11008 11880
rect 10643 11849 10655 11852
rect 10597 11843 10655 11849
rect 9125 11815 9183 11821
rect 9125 11812 9137 11815
rect 8772 11784 9137 11812
rect 8772 11685 8800 11784
rect 9125 11781 9137 11784
rect 9171 11781 9183 11815
rect 9125 11775 9183 11781
rect 9766 11772 9772 11824
rect 9824 11772 9830 11824
rect 10980 11821 11008 11852
rect 11241 11849 11253 11883
rect 11287 11880 11299 11883
rect 12894 11880 12900 11892
rect 11287 11852 12900 11880
rect 11287 11849 11299 11852
rect 11241 11843 11299 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 10965 11815 11023 11821
rect 10965 11781 10977 11815
rect 11011 11781 11023 11815
rect 10965 11775 11023 11781
rect 8527 11648 8708 11676
rect 8757 11679 8815 11685
rect 8527 11645 8539 11648
rect 8481 11639 8539 11645
rect 8757 11645 8769 11679
rect 8803 11645 8815 11679
rect 8757 11639 8815 11645
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 8404 11580 8800 11608
rect 8772 11552 8800 11580
rect 8864 11552 8892 11639
rect 2866 11540 2872 11552
rect 2332 11512 2872 11540
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 3234 11500 3240 11552
rect 3292 11500 3298 11552
rect 3418 11500 3424 11552
rect 3476 11500 3482 11552
rect 5442 11500 5448 11552
rect 5500 11500 5506 11552
rect 5537 11543 5595 11549
rect 5537 11509 5549 11543
rect 5583 11540 5595 11543
rect 5626 11540 5632 11552
rect 5583 11512 5632 11540
rect 5583 11509 5595 11512
rect 5537 11503 5595 11509
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 6638 11500 6644 11552
rect 6696 11500 6702 11552
rect 8754 11500 8760 11552
rect 8812 11500 8818 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9582 11540 9588 11552
rect 8904 11512 9588 11540
rect 8904 11500 8910 11512
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 1104 11450 11868 11472
rect 1104 11398 2295 11450
rect 2347 11398 2359 11450
rect 2411 11398 2423 11450
rect 2475 11398 2487 11450
rect 2539 11398 2551 11450
rect 2603 11398 4986 11450
rect 5038 11398 5050 11450
rect 5102 11398 5114 11450
rect 5166 11398 5178 11450
rect 5230 11398 5242 11450
rect 5294 11398 7677 11450
rect 7729 11398 7741 11450
rect 7793 11398 7805 11450
rect 7857 11398 7869 11450
rect 7921 11398 7933 11450
rect 7985 11398 10368 11450
rect 10420 11398 10432 11450
rect 10484 11398 10496 11450
rect 10548 11398 10560 11450
rect 10612 11398 10624 11450
rect 10676 11398 11868 11450
rect 1104 11376 11868 11398
rect 3234 11296 3240 11348
rect 3292 11296 3298 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4617 11339 4675 11345
rect 4617 11336 4629 11339
rect 4120 11308 4629 11336
rect 4120 11296 4126 11308
rect 4617 11305 4629 11308
rect 4663 11305 4675 11339
rect 4617 11299 4675 11305
rect 5156 11339 5214 11345
rect 5156 11305 5168 11339
rect 5202 11336 5214 11339
rect 5626 11336 5632 11348
rect 5202 11308 5632 11336
rect 5202 11305 5214 11308
rect 5156 11299 5214 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 8662 11336 8668 11348
rect 8527 11308 8668 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 9766 11296 9772 11348
rect 9824 11296 9830 11348
rect 8680 11268 8708 11296
rect 8680 11240 9536 11268
rect 2130 11160 2136 11212
rect 2188 11200 2194 11212
rect 2869 11203 2927 11209
rect 2869 11200 2881 11203
rect 2188 11172 2881 11200
rect 2188 11160 2194 11172
rect 2869 11169 2881 11172
rect 2915 11169 2927 11203
rect 2869 11163 2927 11169
rect 3145 11203 3203 11209
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 4893 11203 4951 11209
rect 4893 11200 4905 11203
rect 3191 11172 4905 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 4893 11169 4905 11172
rect 4939 11200 4951 11203
rect 5534 11200 5540 11212
rect 4939 11172 5540 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 5534 11160 5540 11172
rect 5592 11200 5598 11212
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 5592 11172 6745 11200
rect 5592 11160 5598 11172
rect 6733 11169 6745 11172
rect 6779 11200 6791 11203
rect 8846 11200 8852 11212
rect 6779 11172 8852 11200
rect 6779 11169 6791 11172
rect 6733 11163 6791 11169
rect 8846 11160 8852 11172
rect 8904 11160 8910 11212
rect 9508 11209 9536 11240
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 3513 11135 3571 11141
rect 3513 11132 3525 11135
rect 3160 11104 3525 11132
rect 2406 11024 2412 11076
rect 2464 11024 2470 11076
rect 3160 11064 3188 11104
rect 3513 11101 3525 11104
rect 3559 11101 3571 11135
rect 3513 11095 3571 11101
rect 3602 11092 3608 11144
rect 3660 11132 3666 11144
rect 4341 11135 4399 11141
rect 4341 11132 4353 11135
rect 3660 11104 4353 11132
rect 3660 11092 3666 11104
rect 4341 11101 4353 11104
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 6638 11132 6644 11144
rect 6302 11104 6644 11132
rect 4709 11095 4767 11101
rect 2792 11036 3188 11064
rect 3237 11067 3295 11073
rect 2792 11008 2820 11036
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 4724 11064 4752 11095
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 8757 11135 8815 11141
rect 8757 11132 8769 11135
rect 8352 11104 8769 11132
rect 8352 11092 8358 11104
rect 8757 11101 8769 11104
rect 8803 11101 8815 11135
rect 8757 11095 8815 11101
rect 3283 11036 4660 11064
rect 4724 11036 5488 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 3528 11008 3556 11036
rect 1397 10999 1455 11005
rect 1397 10965 1409 10999
rect 1443 10996 1455 10999
rect 1854 10996 1860 11008
rect 1443 10968 1860 10996
rect 1443 10965 1455 10968
rect 1397 10959 1455 10965
rect 1854 10956 1860 10968
rect 1912 10956 1918 11008
rect 2774 10956 2780 11008
rect 2832 10956 2838 11008
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 3421 10999 3479 11005
rect 3421 10996 3433 10999
rect 3384 10968 3433 10996
rect 3384 10956 3390 10968
rect 3421 10965 3433 10968
rect 3467 10965 3479 10999
rect 3421 10959 3479 10965
rect 3510 10956 3516 11008
rect 3568 10956 3574 11008
rect 3786 10956 3792 11008
rect 3844 10956 3850 11008
rect 4632 10996 4660 11036
rect 5460 11008 5488 11036
rect 7006 11024 7012 11076
rect 7064 11024 7070 11076
rect 8665 11067 8723 11073
rect 8665 11064 8677 11067
rect 8234 11036 8677 11064
rect 8665 11033 8677 11036
rect 8711 11033 8723 11067
rect 8772 11064 8800 11095
rect 9674 11092 9680 11144
rect 9732 11092 9738 11144
rect 10134 11092 10140 11144
rect 10192 11092 10198 11144
rect 9766 11064 9772 11076
rect 8772 11036 9772 11064
rect 8665 11027 8723 11033
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 4706 10996 4712 11008
rect 4632 10968 4712 10996
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 5442 10956 5448 11008
rect 5500 10956 5506 11008
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6641 10999 6699 11005
rect 6641 10996 6653 10999
rect 6052 10968 6653 10996
rect 6052 10956 6058 10968
rect 6641 10965 6653 10968
rect 6687 10965 6699 10999
rect 6641 10959 6699 10965
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 8754 10996 8760 11008
rect 6788 10968 8760 10996
rect 6788 10956 6794 10968
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 8938 10956 8944 11008
rect 8996 10956 9002 11008
rect 9950 10956 9956 11008
rect 10008 10956 10014 11008
rect 1104 10906 11868 10928
rect 1104 10854 2955 10906
rect 3007 10854 3019 10906
rect 3071 10854 3083 10906
rect 3135 10854 3147 10906
rect 3199 10854 3211 10906
rect 3263 10854 5646 10906
rect 5698 10854 5710 10906
rect 5762 10854 5774 10906
rect 5826 10854 5838 10906
rect 5890 10854 5902 10906
rect 5954 10854 8337 10906
rect 8389 10854 8401 10906
rect 8453 10854 8465 10906
rect 8517 10854 8529 10906
rect 8581 10854 8593 10906
rect 8645 10854 11028 10906
rect 11080 10854 11092 10906
rect 11144 10854 11156 10906
rect 11208 10854 11220 10906
rect 11272 10854 11284 10906
rect 11336 10854 11868 10906
rect 1104 10832 11868 10854
rect 2406 10752 2412 10804
rect 2464 10752 2470 10804
rect 3510 10792 3516 10804
rect 2746 10764 3516 10792
rect 2498 10616 2504 10668
rect 2556 10616 2562 10668
rect 2746 10665 2774 10764
rect 3510 10752 3516 10764
rect 3568 10752 3574 10804
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4522 10792 4528 10804
rect 4019 10764 4528 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 5350 10752 5356 10804
rect 5408 10792 5414 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 5408 10764 5457 10792
rect 5408 10752 5414 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 5994 10792 6000 10804
rect 5859 10764 6000 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 6549 10795 6607 10801
rect 6549 10761 6561 10795
rect 6595 10792 6607 10795
rect 6914 10792 6920 10804
rect 6595 10764 6920 10792
rect 6595 10761 6607 10764
rect 6549 10755 6607 10761
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 7064 10764 7113 10792
rect 7064 10752 7070 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 8481 10795 8539 10801
rect 8481 10792 8493 10795
rect 7101 10755 7159 10761
rect 7208 10764 8493 10792
rect 7208 10724 7236 10764
rect 8481 10761 8493 10764
rect 8527 10761 8539 10795
rect 8481 10755 8539 10761
rect 11333 10795 11391 10801
rect 11333 10761 11345 10795
rect 11379 10792 11391 10795
rect 11422 10792 11428 10804
rect 11379 10764 11428 10792
rect 11379 10761 11391 10764
rect 11333 10755 11391 10761
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 7653 10727 7711 10733
rect 7653 10724 7665 10727
rect 3344 10696 4385 10724
rect 3344 10668 3372 10696
rect 2746 10659 2807 10665
rect 2746 10628 2761 10659
rect 2749 10625 2761 10628
rect 2795 10625 2807 10659
rect 2749 10619 2807 10625
rect 3050 10616 3056 10668
rect 3108 10656 3114 10668
rect 3326 10656 3332 10668
rect 3108 10628 3332 10656
rect 3108 10616 3114 10628
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10656 3479 10659
rect 3510 10656 3516 10668
rect 3467 10628 3516 10656
rect 3467 10625 3479 10628
rect 3421 10619 3479 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3602 10616 3608 10668
rect 3660 10616 3666 10668
rect 3694 10616 3700 10668
rect 3752 10616 3758 10668
rect 3786 10616 3792 10668
rect 3844 10616 3850 10668
rect 4357 10665 4385 10696
rect 6656 10696 7236 10724
rect 7300 10696 7665 10724
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 4522 10616 4528 10668
rect 4580 10616 4586 10668
rect 4706 10616 4712 10668
rect 4764 10616 4770 10668
rect 4798 10616 4804 10668
rect 4856 10616 4862 10668
rect 6656 10665 6684 10696
rect 6457 10659 6515 10665
rect 6457 10625 6469 10659
rect 6503 10625 6515 10659
rect 6457 10619 6515 10625
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 6822 10656 6828 10668
rect 6779 10628 6828 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 2915 10591 2973 10597
rect 2915 10588 2927 10591
rect 2792 10560 2927 10588
rect 2792 10532 2820 10560
rect 2915 10557 2927 10560
rect 2961 10557 2973 10591
rect 2915 10551 2973 10557
rect 3142 10548 3148 10600
rect 3200 10548 3206 10600
rect 3712 10588 3740 10616
rect 4154 10588 4160 10600
rect 3712 10560 4160 10588
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10557 4307 10591
rect 4249 10551 4307 10557
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10588 4491 10591
rect 4724 10588 4752 10616
rect 4479 10560 4752 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 2774 10480 2780 10532
rect 2832 10480 2838 10532
rect 3050 10480 3056 10532
rect 3108 10480 3114 10532
rect 3160 10520 3188 10548
rect 4065 10523 4123 10529
rect 4065 10520 4077 10523
rect 3160 10492 4077 10520
rect 4065 10489 4077 10492
rect 4111 10489 4123 10523
rect 4065 10483 4123 10489
rect 2792 10452 2820 10480
rect 4265 10452 4293 10551
rect 5902 10548 5908 10600
rect 5960 10548 5966 10600
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10557 6147 10591
rect 6472 10588 6500 10619
rect 6748 10588 6776 10619
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7300 10656 7328 10696
rect 7653 10693 7665 10696
rect 7699 10693 7711 10727
rect 7653 10687 7711 10693
rect 7745 10727 7803 10733
rect 7745 10693 7757 10727
rect 7791 10724 7803 10727
rect 8938 10724 8944 10736
rect 7791 10696 8944 10724
rect 7791 10693 7803 10696
rect 7745 10687 7803 10693
rect 7009 10619 7067 10625
rect 7116 10628 7328 10656
rect 6472 10560 6776 10588
rect 6089 10551 6147 10557
rect 4338 10480 4344 10532
rect 4396 10520 4402 10532
rect 5077 10523 5135 10529
rect 5077 10520 5089 10523
rect 4396 10492 5089 10520
rect 4396 10480 4402 10492
rect 5077 10489 5089 10492
rect 5123 10520 5135 10523
rect 6104 10520 6132 10551
rect 6638 10520 6644 10532
rect 5123 10492 6644 10520
rect 5123 10489 5135 10492
rect 5077 10483 5135 10489
rect 6638 10480 6644 10492
rect 6696 10480 6702 10532
rect 7024 10520 7052 10619
rect 7116 10600 7144 10628
rect 7374 10616 7380 10668
rect 7432 10616 7438 10668
rect 7668 10656 7696 10687
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 9861 10727 9919 10733
rect 9861 10693 9873 10727
rect 9907 10724 9919 10727
rect 9950 10724 9956 10736
rect 9907 10696 9956 10724
rect 9907 10693 9919 10696
rect 9861 10687 9919 10693
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 10870 10684 10876 10736
rect 10928 10684 10934 10736
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7668 10628 8033 10656
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 7098 10548 7104 10600
rect 7156 10548 7162 10600
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 7300 10520 7328 10551
rect 8220 10532 8248 10619
rect 8294 10616 8300 10668
rect 8352 10616 8358 10668
rect 8386 10616 8392 10668
rect 8444 10616 8450 10668
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10656 8631 10659
rect 8662 10656 8668 10668
rect 8619 10628 8668 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 9582 10548 9588 10600
rect 9640 10548 9646 10600
rect 7837 10523 7895 10529
rect 7837 10520 7849 10523
rect 7024 10492 7144 10520
rect 7300 10492 7849 10520
rect 2792 10424 4293 10452
rect 6730 10412 6736 10464
rect 6788 10412 6794 10464
rect 7116 10452 7144 10492
rect 7837 10489 7849 10492
rect 7883 10489 7895 10523
rect 7837 10483 7895 10489
rect 8202 10480 8208 10532
rect 8260 10480 8266 10532
rect 8294 10452 8300 10464
rect 7116 10424 8300 10452
rect 8294 10412 8300 10424
rect 8352 10452 8358 10464
rect 9490 10452 9496 10464
rect 8352 10424 9496 10452
rect 8352 10412 8358 10424
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 1104 10362 11868 10384
rect 1104 10310 2295 10362
rect 2347 10310 2359 10362
rect 2411 10310 2423 10362
rect 2475 10310 2487 10362
rect 2539 10310 2551 10362
rect 2603 10310 4986 10362
rect 5038 10310 5050 10362
rect 5102 10310 5114 10362
rect 5166 10310 5178 10362
rect 5230 10310 5242 10362
rect 5294 10310 7677 10362
rect 7729 10310 7741 10362
rect 7793 10310 7805 10362
rect 7857 10310 7869 10362
rect 7921 10310 7933 10362
rect 7985 10310 10368 10362
rect 10420 10310 10432 10362
rect 10484 10310 10496 10362
rect 10548 10310 10560 10362
rect 10612 10310 10624 10362
rect 10676 10310 11868 10362
rect 1104 10288 11868 10310
rect 2774 10208 2780 10260
rect 2832 10208 2838 10260
rect 2958 10208 2964 10260
rect 3016 10208 3022 10260
rect 3421 10251 3479 10257
rect 3421 10217 3433 10251
rect 3467 10248 3479 10251
rect 3602 10248 3608 10260
rect 3467 10220 3608 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 3970 10248 3976 10260
rect 3752 10220 3976 10248
rect 3752 10208 3758 10220
rect 3970 10208 3976 10220
rect 4028 10248 4034 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 4028 10220 4169 10248
rect 4028 10208 4034 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 4157 10211 4215 10217
rect 4522 10208 4528 10260
rect 4580 10248 4586 10260
rect 4985 10251 5043 10257
rect 4985 10248 4997 10251
rect 4580 10220 4997 10248
rect 4580 10208 4586 10220
rect 4985 10217 4997 10220
rect 5031 10217 5043 10251
rect 4985 10211 5043 10217
rect 3050 10140 3056 10192
rect 3108 10140 3114 10192
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 3789 10183 3847 10189
rect 3789 10180 3801 10183
rect 3568 10152 3801 10180
rect 3568 10140 3574 10152
rect 3789 10149 3801 10152
rect 3835 10149 3847 10183
rect 5000 10180 5028 10211
rect 5902 10208 5908 10260
rect 5960 10208 5966 10260
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 6880 10220 7205 10248
rect 6880 10208 6886 10220
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 7193 10211 7251 10217
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7432 10220 7665 10248
rect 7432 10208 7438 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 7653 10211 7711 10217
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10229 10251 10287 10257
rect 10229 10248 10241 10251
rect 10192 10220 10241 10248
rect 10192 10208 10198 10220
rect 10229 10217 10241 10220
rect 10275 10217 10287 10251
rect 10229 10211 10287 10217
rect 10870 10208 10876 10260
rect 10928 10208 10934 10260
rect 7098 10180 7104 10192
rect 5000 10152 7104 10180
rect 3789 10143 3847 10149
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 8386 10180 8392 10192
rect 7392 10152 8392 10180
rect 3068 10112 3096 10140
rect 3878 10112 3884 10124
rect 3068 10084 3372 10112
rect 1854 10004 1860 10056
rect 1912 10004 1918 10056
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 2498 10044 2504 10056
rect 2455 10016 2504 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 3344 10053 3372 10084
rect 3528 10084 3884 10112
rect 3528 10053 3556 10084
rect 3878 10072 3884 10084
rect 3936 10112 3942 10124
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 3936 10084 4261 10112
rect 3936 10072 3942 10084
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 4249 10075 4307 10081
rect 5534 10072 5540 10124
rect 5592 10072 5598 10124
rect 6730 10072 6736 10124
rect 6788 10072 6794 10124
rect 2869 10047 2927 10053
rect 2869 10044 2881 10047
rect 2608 10016 2881 10044
rect 1872 9976 1900 10004
rect 2608 9985 2636 10016
rect 2869 10013 2881 10016
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10013 3571 10047
rect 3513 10007 3571 10013
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 4062 10044 4068 10056
rect 4019 10016 4068 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 2593 9979 2651 9985
rect 2593 9976 2605 9979
rect 1872 9948 2605 9976
rect 2593 9945 2605 9948
rect 2639 9945 2651 9979
rect 2593 9939 2651 9945
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 3068 9976 3096 10007
rect 2740 9948 3096 9976
rect 3344 9976 3372 10007
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4798 10044 4804 10056
rect 4264 10016 4804 10044
rect 3694 9976 3700 9988
rect 3344 9948 3700 9976
rect 2740 9936 2746 9948
rect 3694 9936 3700 9948
rect 3752 9936 3758 9988
rect 4264 9920 4292 10016
rect 4798 10004 4804 10016
rect 4856 10044 4862 10056
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4856 10016 4905 10044
rect 4856 10004 4862 10016
rect 4893 10013 4905 10016
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10044 5687 10047
rect 6748 10044 6776 10072
rect 7392 10053 7420 10152
rect 8386 10140 8392 10152
rect 8444 10180 8450 10192
rect 9306 10180 9312 10192
rect 8444 10152 9312 10180
rect 8444 10140 8450 10152
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 9858 10180 9864 10192
rect 9692 10152 9864 10180
rect 8202 10112 8208 10124
rect 7484 10084 8208 10112
rect 5675 10016 6776 10044
rect 7377 10047 7435 10053
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 7377 10013 7389 10047
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 7392 9976 7420 10007
rect 4908 9948 7420 9976
rect 4908 9920 4936 9948
rect 1578 9868 1584 9920
rect 1636 9908 1642 9920
rect 4246 9908 4252 9920
rect 1636 9880 4252 9908
rect 1636 9868 1642 9880
rect 4246 9868 4252 9880
rect 4304 9868 4310 9920
rect 4890 9868 4896 9920
rect 4948 9868 4954 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7484 9908 7512 10084
rect 7852 10053 7880 10084
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8754 10072 8760 10124
rect 8812 10112 8818 10124
rect 9692 10121 9720 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 8812 10084 9689 10112
rect 8812 10072 8818 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 6972 9880 7512 9908
rect 7576 9908 7604 10007
rect 7668 9976 7696 10007
rect 8294 10004 8300 10056
rect 8352 10004 8358 10056
rect 9784 10044 9812 10072
rect 10686 10044 10692 10056
rect 9784 10016 10692 10044
rect 10686 10004 10692 10016
rect 10744 10044 10750 10056
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10744 10016 10977 10044
rect 10744 10004 10750 10016
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 11422 10044 11428 10056
rect 10965 10007 11023 10013
rect 11072 10016 11428 10044
rect 8312 9976 8340 10004
rect 7668 9948 8340 9976
rect 9861 9979 9919 9985
rect 9861 9945 9873 9979
rect 9907 9976 9919 9979
rect 9950 9976 9956 9988
rect 9907 9948 9956 9976
rect 9907 9945 9919 9948
rect 9861 9939 9919 9945
rect 9950 9936 9956 9948
rect 10008 9976 10014 9988
rect 11072 9976 11100 10016
rect 11422 10004 11428 10016
rect 11480 10004 11486 10056
rect 10008 9948 11100 9976
rect 11149 9979 11207 9985
rect 10008 9936 10014 9948
rect 11149 9945 11161 9979
rect 11195 9976 11207 9979
rect 11514 9976 11520 9988
rect 11195 9948 11520 9976
rect 11195 9945 11207 9948
rect 11149 9939 11207 9945
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 8662 9908 8668 9920
rect 7576 9880 8668 9908
rect 6972 9868 6978 9880
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9769 9911 9827 9917
rect 9769 9908 9781 9911
rect 9732 9880 9781 9908
rect 9732 9868 9738 9880
rect 9769 9877 9781 9880
rect 9815 9877 9827 9911
rect 9769 9871 9827 9877
rect 11425 9911 11483 9917
rect 11425 9877 11437 9911
rect 11471 9908 11483 9911
rect 11471 9880 12112 9908
rect 11471 9877 11483 9880
rect 11425 9871 11483 9877
rect 1104 9818 11868 9840
rect 1104 9766 2955 9818
rect 3007 9766 3019 9818
rect 3071 9766 3083 9818
rect 3135 9766 3147 9818
rect 3199 9766 3211 9818
rect 3263 9766 5646 9818
rect 5698 9766 5710 9818
rect 5762 9766 5774 9818
rect 5826 9766 5838 9818
rect 5890 9766 5902 9818
rect 5954 9766 8337 9818
rect 8389 9766 8401 9818
rect 8453 9766 8465 9818
rect 8517 9766 8529 9818
rect 8581 9766 8593 9818
rect 8645 9766 11028 9818
rect 11080 9766 11092 9818
rect 11144 9766 11156 9818
rect 11208 9766 11220 9818
rect 11272 9766 11284 9818
rect 11336 9766 11868 9818
rect 1104 9744 11868 9766
rect 12084 9716 12112 9880
rect 9766 9704 9772 9716
rect 9232 9676 9772 9704
rect 2409 9639 2467 9645
rect 2409 9605 2421 9639
rect 2455 9636 2467 9639
rect 2682 9636 2688 9648
rect 2455 9608 2688 9636
rect 2455 9605 2467 9608
rect 2409 9599 2467 9605
rect 2682 9596 2688 9608
rect 2740 9596 2746 9648
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 7006 9636 7012 9648
rect 5592 9608 7012 9636
rect 5592 9596 5598 9608
rect 7006 9596 7012 9608
rect 7064 9636 7070 9648
rect 9122 9636 9128 9648
rect 7064 9608 9128 9636
rect 7064 9596 7070 9608
rect 9122 9596 9128 9608
rect 9180 9636 9186 9648
rect 9232 9636 9260 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 9950 9664 9956 9716
rect 10008 9664 10014 9716
rect 12066 9664 12072 9716
rect 12124 9664 12130 9716
rect 9180 9608 9260 9636
rect 9180 9596 9186 9608
rect 9306 9596 9312 9648
rect 9364 9596 9370 9648
rect 9493 9639 9551 9645
rect 9493 9605 9505 9639
rect 9539 9636 9551 9639
rect 9968 9636 9996 9664
rect 9539 9608 9996 9636
rect 9539 9605 9551 9608
rect 9493 9599 9551 9605
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 3418 9568 3424 9580
rect 2639 9540 3424 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8772 9540 8861 9568
rect 8772 9376 8800 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 9324 9568 9352 9596
rect 9766 9568 9772 9580
rect 9324 9540 9772 9568
rect 8849 9531 8907 9537
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 9968 9577 9996 9608
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 8938 9460 8944 9512
rect 8996 9460 9002 9512
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9674 9500 9680 9512
rect 9263 9472 9680 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 8904 9404 11560 9432
rect 8904 9392 8910 9404
rect 11532 9376 11560 9404
rect 2777 9367 2835 9373
rect 2777 9333 2789 9367
rect 2823 9364 2835 9367
rect 3602 9364 3608 9376
rect 2823 9336 3608 9364
rect 2823 9333 2835 9336
rect 2777 9327 2835 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 8754 9324 8760 9376
rect 8812 9324 8818 9376
rect 9674 9324 9680 9376
rect 9732 9324 9738 9376
rect 9861 9367 9919 9373
rect 9861 9333 9873 9367
rect 9907 9364 9919 9367
rect 9950 9364 9956 9376
rect 9907 9336 9956 9364
rect 9907 9333 9919 9336
rect 9861 9327 9919 9333
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 11514 9324 11520 9376
rect 11572 9324 11578 9376
rect 1104 9274 11868 9296
rect 1104 9222 2295 9274
rect 2347 9222 2359 9274
rect 2411 9222 2423 9274
rect 2475 9222 2487 9274
rect 2539 9222 2551 9274
rect 2603 9222 4986 9274
rect 5038 9222 5050 9274
rect 5102 9222 5114 9274
rect 5166 9222 5178 9274
rect 5230 9222 5242 9274
rect 5294 9222 7677 9274
rect 7729 9222 7741 9274
rect 7793 9222 7805 9274
rect 7857 9222 7869 9274
rect 7921 9222 7933 9274
rect 7985 9222 10368 9274
rect 10420 9222 10432 9274
rect 10484 9222 10496 9274
rect 10548 9222 10560 9274
rect 10612 9222 10624 9274
rect 10676 9222 11868 9274
rect 1104 9200 11868 9222
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 4154 9160 4160 9172
rect 3283 9132 4160 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 5350 9160 5356 9172
rect 4764 9132 5356 9160
rect 4764 9120 4770 9132
rect 5350 9120 5356 9132
rect 5408 9160 5414 9172
rect 6641 9163 6699 9169
rect 6641 9160 6653 9163
rect 5408 9132 6653 9160
rect 5408 9120 5414 9132
rect 6641 9129 6653 9132
rect 6687 9160 6699 9163
rect 8846 9160 8852 9172
rect 6687 9132 8852 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 9674 9120 9680 9172
rect 9732 9120 9738 9172
rect 10042 9120 10048 9172
rect 10100 9120 10106 9172
rect 3344 8996 3924 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 3344 8965 3372 8996
rect 3896 8968 3924 8996
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 3510 8956 3516 8968
rect 3467 8928 3516 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 2038 8848 2044 8900
rect 2096 8848 2102 8900
rect 2409 8891 2467 8897
rect 2409 8857 2421 8891
rect 2455 8857 2467 8891
rect 3068 8888 3096 8919
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 3620 8888 3648 8919
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3752 8928 3801 8956
rect 3752 8916 3758 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3936 8928 4077 8956
rect 3936 8916 3942 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4172 8956 4200 9120
rect 8665 9095 8723 9101
rect 8665 9061 8677 9095
rect 8711 9092 8723 9095
rect 8938 9092 8944 9104
rect 8711 9064 8944 9092
rect 8711 9061 8723 9064
rect 8665 9055 8723 9061
rect 8938 9052 8944 9064
rect 8996 9092 9002 9104
rect 9398 9092 9404 9104
rect 8996 9064 9404 9092
rect 8996 9052 9002 9064
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 9490 9052 9496 9104
rect 9548 9092 9554 9104
rect 9692 9092 9720 9120
rect 9548 9064 9628 9092
rect 9692 9064 10456 9092
rect 9548 9052 9554 9064
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 9024 4951 9027
rect 6362 9024 6368 9036
rect 4939 8996 6368 9024
rect 4939 8993 4951 8996
rect 4893 8987 4951 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 7006 8984 7012 9036
rect 7064 8984 7070 9036
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 9600 9024 9628 9064
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 8812 8996 9536 9024
rect 9600 8996 9689 9024
rect 8812 8984 8818 8996
rect 4249 8959 4307 8965
rect 4249 8956 4261 8959
rect 4172 8928 4261 8956
rect 4065 8919 4123 8925
rect 4249 8925 4261 8928
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8956 6975 8959
rect 7024 8956 7052 8984
rect 6963 8928 7052 8956
rect 8481 8959 8539 8965
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 8481 8925 8493 8959
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 3068 8860 3648 8888
rect 2409 8851 2467 8857
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 2056 8820 2084 8848
rect 1627 8792 2084 8820
rect 2424 8820 2452 8851
rect 3344 8832 3372 8860
rect 2774 8820 2780 8832
rect 2424 8792 2780 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 2866 8780 2872 8832
rect 2924 8780 2930 8832
rect 3326 8780 3332 8832
rect 3384 8780 3390 8832
rect 3605 8823 3663 8829
rect 3605 8789 3617 8823
rect 3651 8820 3663 8823
rect 3896 8820 3924 8916
rect 4522 8848 4528 8900
rect 4580 8848 4586 8900
rect 4614 8848 4620 8900
rect 4672 8848 4678 8900
rect 5166 8848 5172 8900
rect 5224 8848 5230 8900
rect 6178 8848 6184 8900
rect 6236 8848 6242 8900
rect 8496 8888 8524 8919
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 9324 8965 9352 8996
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8904 8928 8953 8956
rect 8904 8916 8910 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9398 8916 9404 8968
rect 9456 8916 9462 8968
rect 9508 8956 9536 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 9824 8996 9873 9024
rect 9824 8984 9830 8996
rect 9861 8993 9873 8996
rect 9907 8993 9919 9027
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 9861 8987 9919 8993
rect 9968 8996 10333 9024
rect 9968 8956 9996 8996
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 10428 8965 10456 9064
rect 9508 8928 9996 8956
rect 10229 8959 10287 8965
rect 10136 8937 10194 8943
rect 10136 8903 10148 8937
rect 10182 8903 10194 8937
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10136 8900 10194 8903
rect 9769 8891 9827 8897
rect 8496 8860 9628 8888
rect 3651 8792 3924 8820
rect 7009 8823 7067 8829
rect 3651 8789 3663 8792
rect 3605 8783 3663 8789
rect 7009 8789 7021 8823
rect 7055 8820 7067 8823
rect 7098 8820 7104 8832
rect 7055 8792 7104 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 8297 8823 8355 8829
rect 8297 8789 8309 8823
rect 8343 8820 8355 8823
rect 8938 8820 8944 8832
rect 8343 8792 8944 8820
rect 8343 8789 8355 8792
rect 8297 8783 8355 8789
rect 8938 8780 8944 8792
rect 8996 8780 9002 8832
rect 9600 8820 9628 8860
rect 9769 8857 9781 8891
rect 9815 8888 9827 8891
rect 9861 8891 9919 8897
rect 9861 8888 9873 8891
rect 9815 8860 9873 8888
rect 9815 8857 9827 8860
rect 9769 8851 9827 8857
rect 9861 8857 9873 8860
rect 9907 8857 9919 8891
rect 9861 8851 9919 8857
rect 10134 8848 10140 8900
rect 10192 8848 10198 8900
rect 9950 8820 9956 8832
rect 9600 8792 9956 8820
rect 9950 8780 9956 8792
rect 10008 8820 10014 8832
rect 10244 8820 10272 8919
rect 10008 8792 10272 8820
rect 10008 8780 10014 8792
rect 1104 8730 11868 8752
rect 1104 8678 2955 8730
rect 3007 8678 3019 8730
rect 3071 8678 3083 8730
rect 3135 8678 3147 8730
rect 3199 8678 3211 8730
rect 3263 8678 5646 8730
rect 5698 8678 5710 8730
rect 5762 8678 5774 8730
rect 5826 8678 5838 8730
rect 5890 8678 5902 8730
rect 5954 8678 8337 8730
rect 8389 8678 8401 8730
rect 8453 8678 8465 8730
rect 8517 8678 8529 8730
rect 8581 8678 8593 8730
rect 8645 8678 11028 8730
rect 11080 8678 11092 8730
rect 11144 8678 11156 8730
rect 11208 8678 11220 8730
rect 11272 8678 11284 8730
rect 11336 8678 11868 8730
rect 1104 8656 11868 8678
rect 2866 8576 2872 8628
rect 2924 8576 2930 8628
rect 3145 8619 3203 8625
rect 3145 8585 3157 8619
rect 3191 8616 3203 8619
rect 3326 8616 3332 8628
rect 3191 8588 3332 8616
rect 3191 8585 3203 8588
rect 3145 8579 3203 8585
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 4614 8616 4620 8628
rect 3835 8588 4620 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 4706 8576 4712 8628
rect 4764 8576 4770 8628
rect 5166 8576 5172 8628
rect 5224 8576 5230 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6178 8616 6184 8628
rect 6043 8588 6184 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 6472 8588 9628 8616
rect 1762 8440 1768 8492
rect 1820 8480 1826 8492
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1820 8452 2053 8480
rect 1820 8440 1826 8452
rect 2041 8449 2053 8452
rect 2087 8480 2099 8483
rect 2777 8483 2835 8489
rect 2777 8480 2789 8483
rect 2087 8452 2789 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2777 8449 2789 8452
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8412 2191 8415
rect 2884 8412 2912 8576
rect 3418 8548 3424 8560
rect 3068 8520 3424 8548
rect 3068 8489 3096 8520
rect 3418 8508 3424 8520
rect 3476 8548 3482 8560
rect 6472 8548 6500 8588
rect 3476 8520 3648 8548
rect 3476 8508 3482 8520
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 2179 8384 2912 8412
rect 2179 8381 2191 8384
rect 2133 8375 2191 8381
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3252 8412 3280 8443
rect 3510 8440 3516 8492
rect 3568 8440 3574 8492
rect 3620 8489 3648 8520
rect 6380 8520 6500 8548
rect 6380 8492 6408 8520
rect 6546 8508 6552 8560
rect 6604 8548 6610 8560
rect 6641 8551 6699 8557
rect 6641 8548 6653 8551
rect 6604 8520 6653 8548
rect 6604 8508 6610 8520
rect 6641 8517 6653 8520
rect 6687 8517 6699 8551
rect 6641 8511 6699 8517
rect 7098 8508 7104 8560
rect 7156 8508 7162 8560
rect 8665 8551 8723 8557
rect 8665 8517 8677 8551
rect 8711 8548 8723 8551
rect 8846 8548 8852 8560
rect 8711 8520 8852 8548
rect 8711 8517 8723 8520
rect 8665 8511 8723 8517
rect 8846 8508 8852 8520
rect 8904 8508 8910 8560
rect 8938 8508 8944 8560
rect 8996 8508 9002 8560
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8449 3663 8483
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 3605 8443 3663 8449
rect 5092 8452 5365 8480
rect 3789 8415 3847 8421
rect 3789 8412 3801 8415
rect 3016 8384 3801 8412
rect 3016 8372 3022 8384
rect 3789 8381 3801 8384
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 2222 8304 2228 8356
rect 2280 8344 2286 8356
rect 2409 8347 2467 8353
rect 2409 8344 2421 8347
rect 2280 8316 2421 8344
rect 2280 8304 2286 8316
rect 2409 8313 2421 8316
rect 2455 8313 2467 8347
rect 2409 8307 2467 8313
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 3694 8344 3700 8356
rect 2915 8316 3700 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 3694 8304 3700 8316
rect 3752 8304 3758 8356
rect 3804 8288 3832 8375
rect 4246 8372 4252 8424
rect 4304 8412 4310 8424
rect 4433 8415 4491 8421
rect 4433 8412 4445 8415
rect 4304 8384 4445 8412
rect 4304 8372 4310 8384
rect 4433 8381 4445 8384
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 4614 8372 4620 8424
rect 4672 8372 4678 8424
rect 5092 8353 5120 8452
rect 5353 8449 5365 8452
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 5920 8412 5948 8443
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 6086 8412 6092 8424
rect 5920 8384 6092 8412
rect 6086 8372 6092 8384
rect 6144 8412 6150 8424
rect 7006 8412 7012 8424
rect 6144 8384 7012 8412
rect 6144 8372 6150 8384
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8313 5135 8347
rect 5077 8307 5135 8313
rect 8018 8304 8024 8356
rect 8076 8344 8082 8356
rect 8113 8347 8171 8353
rect 8113 8344 8125 8347
rect 8076 8316 8125 8344
rect 8076 8304 8082 8316
rect 8113 8313 8125 8316
rect 8159 8313 8171 8347
rect 8772 8344 8800 8443
rect 8956 8421 8984 8508
rect 9600 8492 9628 8588
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10778 8616 10784 8628
rect 10192 8588 10784 8616
rect 10192 8576 10198 8588
rect 10778 8576 10784 8588
rect 10836 8616 10842 8628
rect 11333 8619 11391 8625
rect 11333 8616 11345 8619
rect 10836 8588 11345 8616
rect 10836 8576 10842 8588
rect 11333 8585 11345 8588
rect 11379 8585 11391 8619
rect 11333 8579 11391 8585
rect 10870 8508 10876 8560
rect 10928 8508 10934 8560
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9582 8440 9588 8492
rect 9640 8440 9646 8492
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 9048 8344 9076 8440
rect 9861 8415 9919 8421
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 10226 8412 10232 8424
rect 9907 8384 10232 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 8772 8316 9076 8344
rect 9401 8347 9459 8353
rect 8113 8307 8171 8313
rect 9401 8313 9413 8347
rect 9447 8344 9459 8347
rect 9447 8316 9720 8344
rect 9447 8313 9459 8316
rect 9401 8307 9459 8313
rect 3786 8236 3792 8288
rect 3844 8236 3850 8288
rect 9692 8276 9720 8316
rect 9858 8276 9864 8288
rect 9692 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 1104 8186 11868 8208
rect 1104 8134 2295 8186
rect 2347 8134 2359 8186
rect 2411 8134 2423 8186
rect 2475 8134 2487 8186
rect 2539 8134 2551 8186
rect 2603 8134 4986 8186
rect 5038 8134 5050 8186
rect 5102 8134 5114 8186
rect 5166 8134 5178 8186
rect 5230 8134 5242 8186
rect 5294 8134 7677 8186
rect 7729 8134 7741 8186
rect 7793 8134 7805 8186
rect 7857 8134 7869 8186
rect 7921 8134 7933 8186
rect 7985 8134 10368 8186
rect 10420 8134 10432 8186
rect 10484 8134 10496 8186
rect 10548 8134 10560 8186
rect 10612 8134 10624 8186
rect 10676 8134 11868 8186
rect 1104 8112 11868 8134
rect 5721 8075 5779 8081
rect 5721 8041 5733 8075
rect 5767 8072 5779 8075
rect 6362 8072 6368 8084
rect 5767 8044 6368 8072
rect 5767 8041 5779 8044
rect 5721 8035 5779 8041
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9030 8072 9036 8084
rect 8987 8044 9036 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 9950 8072 9956 8084
rect 9732 8044 9956 8072
rect 9732 8032 9738 8044
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10226 8032 10232 8084
rect 10284 8072 10290 8084
rect 10413 8075 10471 8081
rect 10413 8072 10425 8075
rect 10284 8044 10425 8072
rect 10284 8032 10290 8044
rect 10413 8041 10425 8044
rect 10459 8041 10471 8075
rect 10413 8035 10471 8041
rect 10870 8032 10876 8084
rect 10928 8032 10934 8084
rect 10321 8007 10379 8013
rect 8312 7976 10088 8004
rect 1946 7896 1952 7948
rect 2004 7936 2010 7948
rect 2317 7939 2375 7945
rect 2317 7936 2329 7939
rect 2004 7908 2329 7936
rect 2004 7896 2010 7908
rect 2317 7905 2329 7908
rect 2363 7936 2375 7939
rect 3510 7936 3516 7948
rect 2363 7908 3516 7936
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 8018 7896 8024 7948
rect 8076 7936 8082 7948
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 8076 7908 8125 7936
rect 8076 7896 8082 7908
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 2038 7828 2044 7880
rect 2096 7828 2102 7880
rect 3418 7828 3424 7880
rect 3476 7828 3482 7880
rect 3602 7828 3608 7880
rect 3660 7828 3666 7880
rect 8312 7877 8340 7976
rect 8662 7896 8668 7948
rect 8720 7936 8726 7948
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 8720 7908 9229 7936
rect 8720 7896 8726 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 9674 7896 9680 7948
rect 9732 7896 9738 7948
rect 9858 7896 9864 7948
rect 9916 7896 9922 7948
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 9122 7868 9128 7880
rect 8619 7840 9128 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 9355 7840 9996 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 1762 7760 1768 7812
rect 1820 7760 1826 7812
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7009 7803 7067 7809
rect 7009 7800 7021 7803
rect 6972 7772 7021 7800
rect 6972 7760 6978 7772
rect 7009 7769 7021 7772
rect 7055 7769 7067 7803
rect 7009 7763 7067 7769
rect 3510 7692 3516 7744
rect 3568 7692 3574 7744
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 9968 7741 9996 7840
rect 10060 7800 10088 7976
rect 10321 7973 10333 8007
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 10336 7868 10364 7967
rect 10686 7964 10692 8016
rect 10744 7964 10750 8016
rect 10597 7871 10655 7877
rect 10597 7868 10609 7871
rect 10336 7840 10609 7868
rect 10597 7837 10609 7840
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 10704 7868 10732 7964
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 10704 7840 10977 7868
rect 10704 7800 10732 7840
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 10060 7772 10732 7800
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7340 7704 7573 7732
rect 7340 7692 7346 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 9953 7735 10011 7741
rect 9953 7701 9965 7735
rect 9999 7732 10011 7735
rect 10778 7732 10784 7744
rect 9999 7704 10784 7732
rect 9999 7701 10011 7704
rect 9953 7695 10011 7701
rect 10778 7692 10784 7704
rect 10836 7692 10842 7744
rect 1104 7642 11868 7664
rect 1104 7590 2955 7642
rect 3007 7590 3019 7642
rect 3071 7590 3083 7642
rect 3135 7590 3147 7642
rect 3199 7590 3211 7642
rect 3263 7590 5646 7642
rect 5698 7590 5710 7642
rect 5762 7590 5774 7642
rect 5826 7590 5838 7642
rect 5890 7590 5902 7642
rect 5954 7590 8337 7642
rect 8389 7590 8401 7642
rect 8453 7590 8465 7642
rect 8517 7590 8529 7642
rect 8581 7590 8593 7642
rect 8645 7590 11028 7642
rect 11080 7590 11092 7642
rect 11144 7590 11156 7642
rect 11208 7590 11220 7642
rect 11272 7590 11284 7642
rect 11336 7590 11868 7642
rect 1104 7568 11868 7590
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 3418 7528 3424 7540
rect 3108 7500 3424 7528
rect 3108 7488 3114 7500
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 3786 7460 3792 7472
rect 3344 7432 3792 7460
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3344 7392 3372 7432
rect 3786 7420 3792 7432
rect 3844 7460 3850 7472
rect 4249 7463 4307 7469
rect 4249 7460 4261 7463
rect 3844 7432 4261 7460
rect 3844 7420 3850 7432
rect 4249 7429 4261 7432
rect 4295 7429 4307 7463
rect 4249 7423 4307 7429
rect 3283 7364 3372 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3344 7336 3372 7364
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3568 7364 3709 7392
rect 3568 7352 3574 7364
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8202 7392 8208 7404
rect 8159 7364 8208 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 3326 7284 3332 7336
rect 3384 7284 3390 7336
rect 3418 7284 3424 7336
rect 3476 7284 3482 7336
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7324 3847 7327
rect 3878 7324 3884 7336
rect 3835 7296 3884 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 4065 7327 4123 7333
rect 4065 7293 4077 7327
rect 4111 7324 4123 7327
rect 4614 7324 4620 7336
rect 4111 7296 4620 7324
rect 4111 7293 4123 7296
rect 4065 7287 4123 7293
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 4212 7160 4537 7188
rect 4212 7148 4218 7160
rect 4525 7157 4537 7160
rect 4571 7188 4583 7191
rect 5534 7188 5540 7200
rect 4571 7160 5540 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 6825 7191 6883 7197
rect 6825 7157 6837 7191
rect 6871 7188 6883 7191
rect 6914 7188 6920 7200
rect 6871 7160 6920 7188
rect 6871 7157 6883 7160
rect 6825 7151 6883 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 1104 7098 11868 7120
rect 1104 7046 2295 7098
rect 2347 7046 2359 7098
rect 2411 7046 2423 7098
rect 2475 7046 2487 7098
rect 2539 7046 2551 7098
rect 2603 7046 4986 7098
rect 5038 7046 5050 7098
rect 5102 7046 5114 7098
rect 5166 7046 5178 7098
rect 5230 7046 5242 7098
rect 5294 7046 7677 7098
rect 7729 7046 7741 7098
rect 7793 7046 7805 7098
rect 7857 7046 7869 7098
rect 7921 7046 7933 7098
rect 7985 7046 10368 7098
rect 10420 7046 10432 7098
rect 10484 7046 10496 7098
rect 10548 7046 10560 7098
rect 10612 7046 10624 7098
rect 10676 7046 11868 7098
rect 1104 7024 11868 7046
rect 3602 6944 3608 6996
rect 3660 6944 3666 6996
rect 6822 6944 6828 6996
rect 6880 6984 6886 6996
rect 7101 6987 7159 6993
rect 7101 6984 7113 6987
rect 6880 6956 7113 6984
rect 6880 6944 6886 6956
rect 7101 6953 7113 6956
rect 7147 6953 7159 6987
rect 7101 6947 7159 6953
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6953 7343 6987
rect 7285 6947 7343 6953
rect 7653 6987 7711 6993
rect 7653 6953 7665 6987
rect 7699 6953 7711 6987
rect 7653 6947 7711 6953
rect 3418 6876 3424 6928
rect 3476 6916 3482 6928
rect 7300 6916 7328 6947
rect 7668 6916 7696 6947
rect 9674 6916 9680 6928
rect 3476 6888 4016 6916
rect 3476 6876 3482 6888
rect 1854 6808 1860 6860
rect 1912 6808 1918 6860
rect 2038 6808 2044 6860
rect 2096 6848 2102 6860
rect 2133 6851 2191 6857
rect 2133 6848 2145 6851
rect 2096 6820 2145 6848
rect 2096 6808 2102 6820
rect 2133 6817 2145 6820
rect 2179 6817 2191 6851
rect 3988 6848 4016 6888
rect 6472 6888 7328 6916
rect 7576 6888 7696 6916
rect 8220 6888 9680 6916
rect 6472 6848 6500 6888
rect 2133 6811 2191 6817
rect 3344 6820 3924 6848
rect 3988 6820 5396 6848
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 1765 6783 1823 6789
rect 1765 6780 1777 6783
rect 1728 6752 1777 6780
rect 1728 6740 1734 6752
rect 1765 6749 1777 6752
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 3050 6740 3056 6792
rect 3108 6740 3114 6792
rect 3344 6789 3372 6820
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3418 6740 3424 6792
rect 3476 6740 3482 6792
rect 3510 6740 3516 6792
rect 3568 6740 3574 6792
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 3237 6715 3295 6721
rect 3237 6681 3249 6715
rect 3283 6712 3295 6715
rect 3528 6712 3556 6740
rect 3283 6684 3556 6712
rect 3283 6681 3295 6684
rect 3237 6675 3295 6681
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 3151 6647 3209 6653
rect 3151 6644 3163 6647
rect 2280 6616 3163 6644
rect 2280 6604 2286 6616
rect 3151 6613 3163 6616
rect 3197 6613 3209 6647
rect 3151 6607 3209 6613
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 3620 6644 3648 6743
rect 3896 6724 3924 6820
rect 5368 6792 5396 6820
rect 5736 6820 6500 6848
rect 6549 6851 6607 6857
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 3878 6672 3884 6724
rect 3936 6672 3942 6724
rect 5166 6672 5172 6724
rect 5224 6712 5230 6724
rect 5736 6712 5764 6820
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7576 6848 7604 6888
rect 8220 6848 8248 6888
rect 9674 6876 9680 6888
rect 9732 6916 9738 6928
rect 9732 6888 10088 6916
rect 9732 6876 9738 6888
rect 6595 6820 7604 6848
rect 7668 6820 8248 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 6089 6783 6147 6789
rect 5859 6752 6040 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 5224 6684 5917 6712
rect 5224 6672 5230 6684
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 5905 6675 5963 6681
rect 6012 6656 6040 6752
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 6822 6780 6828 6792
rect 6687 6752 6828 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 6104 6712 6132 6743
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7282 6780 7288 6792
rect 7055 6752 7288 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7432 6752 7573 6780
rect 7432 6740 7438 6752
rect 7561 6749 7573 6752
rect 7607 6780 7619 6783
rect 7668 6780 7696 6820
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 10060 6857 10088 6888
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9640 6820 9965 6848
rect 9640 6808 9646 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 9953 6811 10011 6817
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 7607 6752 7696 6780
rect 7745 6783 7803 6789
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 7791 6752 8493 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 8481 6749 8493 6752
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8665 6783 8723 6789
rect 8665 6749 8677 6783
rect 8711 6780 8723 6783
rect 8754 6780 8760 6792
rect 8711 6752 8760 6780
rect 8711 6749 8723 6752
rect 8665 6743 8723 6749
rect 7466 6712 7472 6724
rect 6104 6684 7472 6712
rect 7466 6672 7472 6684
rect 7524 6672 7530 6724
rect 7760 6712 7788 6743
rect 7576 6684 7788 6712
rect 8496 6712 8524 6743
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 8956 6712 8984 6743
rect 9122 6740 9128 6792
rect 9180 6740 9186 6792
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9272 6752 9413 6780
rect 9272 6740 9278 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9858 6740 9864 6792
rect 9916 6740 9922 6792
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 8496 6684 8984 6712
rect 7576 6656 7604 6684
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 10152 6712 10180 6743
rect 9548 6684 10180 6712
rect 9548 6672 9554 6684
rect 3384 6616 3648 6644
rect 3384 6604 3390 6616
rect 5994 6604 6000 6656
rect 6052 6604 6058 6656
rect 6270 6604 6276 6656
rect 6328 6604 6334 6656
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6644 6423 6647
rect 6546 6644 6552 6656
rect 6411 6616 6552 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 7282 6653 7288 6656
rect 7269 6647 7288 6653
rect 7269 6613 7281 6647
rect 7269 6607 7288 6613
rect 7282 6604 7288 6607
rect 7340 6604 7346 6656
rect 7558 6604 7564 6656
rect 7616 6604 7622 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 8846 6644 8852 6656
rect 8619 6616 8852 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 9585 6647 9643 6653
rect 9585 6644 9597 6647
rect 9456 6616 9597 6644
rect 9456 6604 9462 6616
rect 9585 6613 9597 6616
rect 9631 6613 9643 6647
rect 9585 6607 9643 6613
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 1104 6554 11868 6576
rect 1104 6502 2955 6554
rect 3007 6502 3019 6554
rect 3071 6502 3083 6554
rect 3135 6502 3147 6554
rect 3199 6502 3211 6554
rect 3263 6502 5646 6554
rect 5698 6502 5710 6554
rect 5762 6502 5774 6554
rect 5826 6502 5838 6554
rect 5890 6502 5902 6554
rect 5954 6502 8337 6554
rect 8389 6502 8401 6554
rect 8453 6502 8465 6554
rect 8517 6502 8529 6554
rect 8581 6502 8593 6554
rect 8645 6502 11028 6554
rect 11080 6502 11092 6554
rect 11144 6502 11156 6554
rect 11208 6502 11220 6554
rect 11272 6502 11284 6554
rect 11336 6502 11868 6554
rect 1104 6480 11868 6502
rect 2222 6400 2228 6452
rect 2280 6400 2286 6452
rect 3329 6443 3387 6449
rect 3329 6409 3341 6443
rect 3375 6440 3387 6443
rect 3510 6440 3516 6452
rect 3375 6412 3516 6440
rect 3375 6409 3387 6412
rect 3329 6403 3387 6409
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 3878 6400 3884 6452
rect 3936 6400 3942 6452
rect 4522 6400 4528 6452
rect 4580 6400 4586 6452
rect 5074 6440 5080 6452
rect 4908 6412 5080 6440
rect 2038 6264 2044 6316
rect 2096 6304 2102 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 2096 6276 2145 6304
rect 2096 6264 2102 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2148 6100 2176 6267
rect 2240 6245 2268 6400
rect 4430 6372 4436 6384
rect 4172 6344 4436 6372
rect 4172 6313 4200 6344
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 4540 6372 4568 6400
rect 4908 6381 4936 6412
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5166 6400 5172 6452
rect 5224 6400 5230 6452
rect 5813 6443 5871 6449
rect 5813 6409 5825 6443
rect 5859 6440 5871 6443
rect 5994 6440 6000 6452
rect 5859 6412 6000 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 5994 6400 6000 6412
rect 6052 6440 6058 6452
rect 7006 6440 7012 6452
rect 6052 6412 7012 6440
rect 6052 6400 6058 6412
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 7147 6412 7504 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 4893 6375 4951 6381
rect 4540 6344 4844 6372
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4338 6264 4344 6316
rect 4396 6304 4402 6316
rect 4540 6313 4568 6344
rect 4816 6313 4844 6344
rect 4893 6341 4905 6375
rect 4939 6341 4951 6375
rect 4893 6335 4951 6341
rect 6270 6332 6276 6384
rect 6328 6372 6334 6384
rect 6733 6375 6791 6381
rect 6733 6372 6745 6375
rect 6328 6344 6500 6372
rect 6328 6332 6334 6344
rect 4518 6307 4576 6313
rect 4396 6276 4476 6304
rect 4396 6264 4402 6276
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6205 2283 6239
rect 2225 6199 2283 6205
rect 3878 6196 3884 6248
rect 3936 6196 3942 6248
rect 4448 6236 4476 6276
rect 4518 6273 4530 6307
rect 4564 6273 4576 6307
rect 4518 6267 4576 6273
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 4847 6276 5089 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 5077 6273 5089 6276
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 4632 6236 4660 6267
rect 5184 6236 5212 6267
rect 5258 6264 5264 6316
rect 5316 6264 5322 6316
rect 5350 6264 5356 6316
rect 5408 6264 5414 6316
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6472 6313 6500 6344
rect 6564 6344 6745 6372
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5592 6276 5825 6304
rect 5592 6264 5598 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6457 6307 6515 6313
rect 6457 6273 6469 6307
rect 6503 6273 6515 6307
rect 6457 6267 6515 6273
rect 4448 6208 5212 6236
rect 2501 6171 2559 6177
rect 2501 6137 2513 6171
rect 2547 6168 2559 6171
rect 2682 6168 2688 6180
rect 2547 6140 2688 6168
rect 2547 6137 2559 6140
rect 2501 6131 2559 6137
rect 2682 6128 2688 6140
rect 2740 6128 2746 6180
rect 2958 6128 2964 6180
rect 3016 6168 3022 6180
rect 4065 6171 4123 6177
rect 4065 6168 4077 6171
rect 3016 6140 4077 6168
rect 3016 6128 3022 6140
rect 4065 6137 4077 6140
rect 4111 6137 4123 6171
rect 5074 6168 5080 6180
rect 4065 6131 4123 6137
rect 4356 6140 5080 6168
rect 3329 6103 3387 6109
rect 3329 6100 3341 6103
rect 2148 6072 3341 6100
rect 3329 6069 3341 6072
rect 3375 6069 3387 6103
rect 3329 6063 3387 6069
rect 3513 6103 3571 6109
rect 3513 6069 3525 6103
rect 3559 6100 3571 6103
rect 4356 6100 4384 6140
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 5368 6168 5396 6264
rect 5828 6236 5856 6267
rect 6564 6236 6592 6344
rect 6733 6341 6745 6344
rect 6779 6372 6791 6375
rect 7476 6372 7504 6412
rect 7558 6400 7564 6452
rect 7616 6400 7622 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8938 6440 8944 6452
rect 8343 6412 8944 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9401 6443 9459 6449
rect 9401 6409 9413 6443
rect 9447 6440 9459 6443
rect 9490 6440 9496 6452
rect 9447 6412 9496 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 9732 6412 9812 6440
rect 9732 6400 9738 6412
rect 8478 6372 8484 6384
rect 6779 6344 7312 6372
rect 7476 6344 7696 6372
rect 6779 6341 6791 6344
rect 6733 6335 6791 6341
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 5828 6208 6592 6236
rect 5426 6171 5484 6177
rect 5426 6168 5438 6171
rect 5368 6140 5438 6168
rect 5426 6137 5438 6140
rect 5472 6137 5484 6171
rect 6656 6168 6684 6267
rect 6748 6236 6776 6335
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6963 6276 7205 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7284 6307 7312 6344
rect 7668 6313 7696 6344
rect 8128 6344 8484 6372
rect 7377 6307 7435 6313
rect 7284 6302 7328 6307
rect 7377 6302 7389 6307
rect 7284 6279 7389 6302
rect 7300 6274 7389 6279
rect 7193 6267 7251 6273
rect 7377 6273 7389 6274
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7477 6305 7535 6311
rect 7477 6271 7489 6305
rect 7523 6302 7535 6305
rect 7653 6307 7711 6313
rect 7523 6274 7604 6302
rect 7523 6271 7535 6274
rect 6822 6236 6828 6248
rect 6748 6208 6828 6236
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7208 6236 7236 6267
rect 7477 6265 7535 6271
rect 7156 6208 7236 6236
rect 7285 6239 7343 6245
rect 7156 6196 7162 6208
rect 7285 6205 7297 6239
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 7300 6168 7328 6199
rect 7576 6168 7604 6274
rect 7653 6273 7665 6307
rect 7699 6273 7711 6307
rect 7653 6267 7711 6273
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8018 6304 8024 6316
rect 7975 6276 8024 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8128 6313 8156 6344
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 9784 6381 9812 6412
rect 9769 6375 9827 6381
rect 9769 6341 9781 6375
rect 9815 6341 9827 6375
rect 9769 6335 9827 6341
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 8294 6264 8300 6316
rect 8352 6304 8358 6316
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8352 6276 8585 6304
rect 8352 6264 8358 6276
rect 8573 6273 8585 6276
rect 8619 6304 8631 6307
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 8619 6276 9229 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 9217 6273 9229 6276
rect 9263 6304 9275 6307
rect 9306 6304 9312 6316
rect 9263 6276 9312 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 10870 6264 10876 6316
rect 10928 6264 10934 6316
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8202 6236 8208 6248
rect 7883 6208 8208 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 8662 6196 8668 6248
rect 8720 6196 8726 6248
rect 9030 6196 9036 6248
rect 9088 6196 9094 6248
rect 9490 6196 9496 6248
rect 9548 6196 9554 6248
rect 9766 6236 9772 6248
rect 9600 6208 9772 6236
rect 9600 6168 9628 6208
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 6656 6140 7604 6168
rect 8864 6140 9628 6168
rect 5426 6131 5484 6137
rect 3559 6072 4384 6100
rect 3559 6069 3571 6072
rect 3513 6063 3571 6069
rect 4430 6060 4436 6112
rect 4488 6060 4494 6112
rect 4798 6060 4804 6112
rect 4856 6060 4862 6112
rect 5534 6060 5540 6112
rect 5592 6060 5598 6112
rect 5626 6060 5632 6112
rect 5684 6060 5690 6112
rect 6549 6103 6607 6109
rect 6549 6069 6561 6103
rect 6595 6100 6607 6103
rect 7006 6100 7012 6112
rect 6595 6072 7012 6100
rect 6595 6069 6607 6072
rect 6549 6063 6607 6069
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 8864 6100 8892 6140
rect 8536 6072 8892 6100
rect 8941 6103 8999 6109
rect 8536 6060 8542 6072
rect 8941 6069 8953 6103
rect 8987 6100 8999 6103
rect 9030 6100 9036 6112
rect 8987 6072 9036 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 9306 6060 9312 6112
rect 9364 6100 9370 6112
rect 11241 6103 11299 6109
rect 11241 6100 11253 6103
rect 9364 6072 11253 6100
rect 9364 6060 9370 6072
rect 11241 6069 11253 6072
rect 11287 6069 11299 6103
rect 11241 6063 11299 6069
rect 1104 6010 11868 6032
rect 1104 5958 2295 6010
rect 2347 5958 2359 6010
rect 2411 5958 2423 6010
rect 2475 5958 2487 6010
rect 2539 5958 2551 6010
rect 2603 5958 4986 6010
rect 5038 5958 5050 6010
rect 5102 5958 5114 6010
rect 5166 5958 5178 6010
rect 5230 5958 5242 6010
rect 5294 5958 7677 6010
rect 7729 5958 7741 6010
rect 7793 5958 7805 6010
rect 7857 5958 7869 6010
rect 7921 5958 7933 6010
rect 7985 5958 10368 6010
rect 10420 5958 10432 6010
rect 10484 5958 10496 6010
rect 10548 5958 10560 6010
rect 10612 5958 10624 6010
rect 10676 5958 11868 6010
rect 1104 5936 11868 5958
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 3878 5856 3884 5908
rect 3936 5856 3942 5908
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4396 5868 4445 5896
rect 4396 5856 4402 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 5074 5896 5080 5908
rect 4764 5868 5080 5896
rect 4764 5856 4770 5868
rect 5074 5856 5080 5868
rect 5132 5896 5138 5908
rect 6914 5896 6920 5908
rect 5132 5868 6920 5896
rect 5132 5856 5138 5868
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 8205 5899 8263 5905
rect 8205 5896 8217 5899
rect 8168 5868 8217 5896
rect 8168 5856 8174 5868
rect 8205 5865 8217 5868
rect 8251 5865 8263 5899
rect 8205 5859 8263 5865
rect 8662 5856 8668 5908
rect 8720 5856 8726 5908
rect 8938 5856 8944 5908
rect 8996 5856 9002 5908
rect 9214 5856 9220 5908
rect 9272 5856 9278 5908
rect 9309 5899 9367 5905
rect 9309 5865 9321 5899
rect 9355 5896 9367 5899
rect 9858 5896 9864 5908
rect 9355 5868 9864 5896
rect 9355 5865 9367 5868
rect 9309 5859 9367 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10686 5856 10692 5908
rect 10744 5856 10750 5908
rect 10870 5856 10876 5908
rect 10928 5856 10934 5908
rect 1872 5760 1900 5856
rect 1949 5763 2007 5769
rect 1949 5760 1961 5763
rect 1872 5732 1961 5760
rect 1949 5729 1961 5732
rect 1995 5760 2007 5763
rect 3326 5760 3332 5772
rect 1995 5732 3332 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2590 5692 2596 5704
rect 2271 5664 2596 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 3896 5624 3924 5856
rect 4080 5800 5488 5828
rect 4080 5701 4108 5800
rect 4154 5720 4160 5772
rect 4212 5720 4218 5772
rect 4890 5720 4896 5772
rect 4948 5760 4954 5772
rect 5460 5769 5488 5800
rect 6822 5788 6828 5840
rect 6880 5828 6886 5840
rect 8680 5828 8708 5856
rect 6880 5800 8708 5828
rect 6880 5788 6886 5800
rect 5261 5763 5319 5769
rect 5261 5760 5273 5763
rect 4948 5732 5273 5760
rect 4948 5720 4954 5732
rect 5261 5729 5273 5732
rect 5307 5729 5319 5763
rect 5261 5723 5319 5729
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5626 5760 5632 5772
rect 5491 5732 5632 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 5626 5720 5632 5732
rect 5684 5760 5690 5772
rect 8570 5760 8576 5772
rect 5684 5732 6316 5760
rect 5684 5720 5690 5732
rect 6288 5704 6316 5732
rect 8036 5732 8576 5760
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 4798 5652 4804 5704
rect 4856 5652 4862 5704
rect 5074 5652 5080 5704
rect 5132 5652 5138 5704
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 8036 5701 8064 5732
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 8297 5695 8355 5701
rect 8297 5692 8309 5695
rect 8260 5664 8309 5692
rect 8260 5652 8266 5664
rect 8297 5661 8309 5664
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8680 5692 8708 5800
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 9232 5828 9260 5856
rect 10704 5828 10732 5856
rect 11149 5831 11207 5837
rect 11149 5828 11161 5831
rect 8803 5800 9260 5828
rect 9324 5800 9812 5828
rect 10704 5800 11161 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 9324 5772 9352 5800
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 8904 5732 8984 5760
rect 8904 5720 8910 5732
rect 8956 5701 8984 5732
rect 9030 5720 9036 5772
rect 9088 5720 9094 5772
rect 9306 5720 9312 5772
rect 9364 5720 9370 5772
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5760 9459 5763
rect 9582 5760 9588 5772
rect 9447 5732 9588 5760
rect 9447 5729 9459 5732
rect 9401 5723 9459 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 9784 5769 9812 5800
rect 9769 5763 9827 5769
rect 9769 5729 9781 5763
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 8527 5664 8708 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 5169 5627 5227 5633
rect 3896 5596 4660 5624
rect 2869 5559 2927 5565
rect 2869 5525 2881 5559
rect 2915 5556 2927 5559
rect 2958 5556 2964 5568
rect 2915 5528 2964 5556
rect 2915 5525 2927 5528
rect 2869 5519 2927 5525
rect 2958 5516 2964 5528
rect 3016 5556 3022 5568
rect 3694 5556 3700 5568
rect 3016 5528 3700 5556
rect 3016 5516 3022 5528
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 4522 5516 4528 5568
rect 4580 5516 4586 5568
rect 4632 5556 4660 5596
rect 5169 5593 5181 5627
rect 5215 5624 5227 5627
rect 5215 5596 5580 5624
rect 5215 5593 5227 5596
rect 5169 5587 5227 5593
rect 5552 5568 5580 5596
rect 7098 5584 7104 5636
rect 7156 5624 7162 5636
rect 8128 5624 8156 5652
rect 8404 5624 8432 5655
rect 7156 5596 8432 5624
rect 8680 5624 8708 5664
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5692 8999 5695
rect 9490 5692 9496 5704
rect 8987 5664 9496 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 10980 5701 11008 5800
rect 11149 5797 11161 5800
rect 11195 5797 11207 5831
rect 11149 5791 11207 5797
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5692 11483 5695
rect 11790 5692 11796 5704
rect 11471 5664 11796 5692
rect 11471 5661 11483 5664
rect 11425 5655 11483 5661
rect 8846 5624 8852 5636
rect 8680 5596 8852 5624
rect 7156 5584 7162 5596
rect 8846 5584 8852 5596
rect 8904 5584 8910 5636
rect 9766 5584 9772 5636
rect 9824 5624 9830 5636
rect 9876 5624 9904 5655
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 9824 5596 9904 5624
rect 9824 5584 9830 5596
rect 5261 5559 5319 5565
rect 5261 5556 5273 5559
rect 4632 5528 5273 5556
rect 5261 5525 5273 5528
rect 5307 5525 5319 5559
rect 5261 5519 5319 5525
rect 5534 5516 5540 5568
rect 5592 5516 5598 5568
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 9398 5556 9404 5568
rect 8996 5528 9404 5556
rect 8996 5516 9002 5528
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 10042 5516 10048 5568
rect 10100 5516 10106 5568
rect 1104 5466 11868 5488
rect 1104 5414 2955 5466
rect 3007 5414 3019 5466
rect 3071 5414 3083 5466
rect 3135 5414 3147 5466
rect 3199 5414 3211 5466
rect 3263 5414 5646 5466
rect 5698 5414 5710 5466
rect 5762 5414 5774 5466
rect 5826 5414 5838 5466
rect 5890 5414 5902 5466
rect 5954 5414 8337 5466
rect 8389 5414 8401 5466
rect 8453 5414 8465 5466
rect 8517 5414 8529 5466
rect 8581 5414 8593 5466
rect 8645 5414 11028 5466
rect 11080 5414 11092 5466
rect 11144 5414 11156 5466
rect 11208 5414 11220 5466
rect 11272 5414 11284 5466
rect 11336 5414 11868 5466
rect 1104 5392 11868 5414
rect 2409 5355 2467 5361
rect 2409 5321 2421 5355
rect 2455 5352 2467 5355
rect 2682 5352 2688 5364
rect 2455 5324 2688 5352
rect 2455 5321 2467 5324
rect 2409 5315 2467 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 4706 5312 4712 5364
rect 4764 5312 4770 5364
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 4948 5324 6561 5352
rect 4948 5312 4954 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 9122 5352 9128 5364
rect 8803 5324 9128 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 9398 5312 9404 5364
rect 9456 5312 9462 5364
rect 934 5244 940 5296
rect 992 5284 998 5296
rect 1397 5287 1455 5293
rect 1397 5284 1409 5287
rect 992 5256 1409 5284
rect 992 5244 998 5256
rect 1397 5253 1409 5256
rect 1443 5253 1455 5287
rect 1397 5247 1455 5253
rect 1670 5244 1676 5296
rect 1728 5284 1734 5296
rect 1765 5287 1823 5293
rect 1765 5284 1777 5287
rect 1728 5256 1777 5284
rect 1728 5244 1734 5256
rect 1765 5253 1777 5256
rect 1811 5284 1823 5287
rect 2317 5287 2375 5293
rect 2317 5284 2329 5287
rect 1811 5256 2329 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 2317 5253 2329 5256
rect 2363 5284 2375 5287
rect 3326 5284 3332 5296
rect 2363 5256 3332 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 3326 5244 3332 5256
rect 3384 5284 3390 5296
rect 3384 5256 4660 5284
rect 3384 5244 3390 5256
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 2096 5120 2513 5148
rect 2096 5108 2102 5120
rect 2501 5117 2513 5120
rect 2547 5148 2559 5151
rect 2547 5120 2774 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 1946 4972 1952 5024
rect 2004 4972 2010 5024
rect 2746 5012 2774 5120
rect 4430 5108 4436 5160
rect 4488 5148 4494 5160
rect 4540 5148 4568 5179
rect 4488 5120 4568 5148
rect 4632 5148 4660 5256
rect 4724 5256 7328 5284
rect 4724 5225 4752 5256
rect 7300 5228 7328 5256
rect 9030 5244 9036 5296
rect 9088 5244 9094 5296
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 5350 5176 5356 5228
rect 5408 5176 5414 5228
rect 6457 5219 6515 5225
rect 6457 5185 6469 5219
rect 6503 5216 6515 5219
rect 6822 5216 6828 5228
rect 6503 5188 6828 5216
rect 6503 5185 6515 5188
rect 6457 5179 6515 5185
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 7282 5176 7288 5228
rect 7340 5176 7346 5228
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8812 5188 8953 5216
rect 8812 5176 8818 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 9048 5216 9076 5244
rect 9416 5225 9444 5312
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 9048 5188 9321 5216
rect 8941 5179 8999 5185
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 5368 5148 5396 5176
rect 4632 5120 5396 5148
rect 9324 5148 9352 5179
rect 9490 5176 9496 5228
rect 9548 5176 9554 5228
rect 9677 5151 9735 5157
rect 9677 5148 9689 5151
rect 9324 5120 9689 5148
rect 4488 5108 4494 5120
rect 9677 5117 9689 5120
rect 9723 5117 9735 5151
rect 9677 5111 9735 5117
rect 9582 5040 9588 5092
rect 9640 5040 9646 5092
rect 2866 5012 2872 5024
rect 2746 4984 2872 5012
rect 2866 4972 2872 4984
rect 2924 4972 2930 5024
rect 9214 4972 9220 5024
rect 9272 4972 9278 5024
rect 1104 4922 11868 4944
rect 1104 4870 2295 4922
rect 2347 4870 2359 4922
rect 2411 4870 2423 4922
rect 2475 4870 2487 4922
rect 2539 4870 2551 4922
rect 2603 4870 4986 4922
rect 5038 4870 5050 4922
rect 5102 4870 5114 4922
rect 5166 4870 5178 4922
rect 5230 4870 5242 4922
rect 5294 4870 7677 4922
rect 7729 4870 7741 4922
rect 7793 4870 7805 4922
rect 7857 4870 7869 4922
rect 7921 4870 7933 4922
rect 7985 4870 10368 4922
rect 10420 4870 10432 4922
rect 10484 4870 10496 4922
rect 10548 4870 10560 4922
rect 10612 4870 10624 4922
rect 10676 4870 11868 4922
rect 1104 4848 11868 4870
rect 1946 4768 1952 4820
rect 2004 4768 2010 4820
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5629 4811 5687 4817
rect 5629 4808 5641 4811
rect 5592 4780 5641 4808
rect 5592 4768 5598 4780
rect 5629 4777 5641 4780
rect 5675 4777 5687 4811
rect 5629 4771 5687 4777
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9272 4780 9413 4808
rect 9272 4768 9278 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 1964 4604 1992 4768
rect 7098 4700 7104 4752
rect 7156 4700 7162 4752
rect 7469 4743 7527 4749
rect 7469 4709 7481 4743
rect 7515 4740 7527 4743
rect 8754 4740 8760 4752
rect 7515 4712 8760 4740
rect 7515 4709 7527 4712
rect 7469 4703 7527 4709
rect 4430 4632 4436 4684
rect 4488 4632 4494 4684
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6880 4644 7021 4672
rect 6880 4632 6886 4644
rect 7009 4641 7021 4644
rect 7055 4641 7067 4675
rect 7116 4672 7144 4700
rect 7837 4675 7895 4681
rect 7837 4672 7849 4675
rect 7116 4644 7849 4672
rect 7009 4635 7067 4641
rect 7837 4641 7849 4644
rect 7883 4641 7895 4675
rect 7837 4635 7895 4641
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 1964 4576 2145 4604
rect 2133 4573 2145 4576
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 4890 4564 4896 4616
rect 4948 4564 4954 4616
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 7944 4613 7972 4712
rect 8754 4700 8760 4712
rect 8812 4700 8818 4752
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8904 4644 9045 4672
rect 8904 4632 8910 4644
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 7929 4607 7987 4613
rect 7147 4576 7236 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 4801 4539 4859 4545
rect 4801 4505 4813 4539
rect 4847 4536 4859 4539
rect 6288 4536 6316 4564
rect 4847 4508 6316 4536
rect 4847 4505 4859 4508
rect 4801 4499 4859 4505
rect 7208 4480 7236 4576
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8662 4564 8668 4616
rect 8720 4604 8726 4616
rect 9122 4604 9128 4616
rect 8720 4576 9128 4604
rect 8720 4564 8726 4576
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 9416 4604 9444 4771
rect 10042 4632 10048 4684
rect 10100 4632 10106 4684
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 9416 4576 9965 4604
rect 9953 4573 9965 4576
rect 9999 4573 10011 4607
rect 9953 4567 10011 4573
rect 1946 4428 1952 4480
rect 2004 4428 2010 4480
rect 3786 4428 3792 4480
rect 3844 4468 3850 4480
rect 4709 4471 4767 4477
rect 4709 4468 4721 4471
rect 3844 4440 4721 4468
rect 3844 4428 3850 4440
rect 4709 4437 4721 4440
rect 4755 4437 4767 4471
rect 4709 4431 4767 4437
rect 7190 4428 7196 4480
rect 7248 4428 7254 4480
rect 7558 4428 7564 4480
rect 7616 4428 7622 4480
rect 9582 4428 9588 4480
rect 9640 4428 9646 4480
rect 1104 4378 11868 4400
rect 1104 4326 2955 4378
rect 3007 4326 3019 4378
rect 3071 4326 3083 4378
rect 3135 4326 3147 4378
rect 3199 4326 3211 4378
rect 3263 4326 5646 4378
rect 5698 4326 5710 4378
rect 5762 4326 5774 4378
rect 5826 4326 5838 4378
rect 5890 4326 5902 4378
rect 5954 4326 8337 4378
rect 8389 4326 8401 4378
rect 8453 4326 8465 4378
rect 8517 4326 8529 4378
rect 8581 4326 8593 4378
rect 8645 4326 11028 4378
rect 11080 4326 11092 4378
rect 11144 4326 11156 4378
rect 11208 4326 11220 4378
rect 11272 4326 11284 4378
rect 11336 4326 11868 4378
rect 1104 4304 11868 4326
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 4154 4264 4160 4276
rect 2740 4236 4160 4264
rect 2740 4224 2746 4236
rect 4154 4224 4160 4236
rect 4212 4264 4218 4276
rect 4525 4267 4583 4273
rect 4525 4264 4537 4267
rect 4212 4236 4537 4264
rect 4212 4224 4218 4236
rect 4525 4233 4537 4236
rect 4571 4264 4583 4267
rect 5442 4264 5448 4276
rect 4571 4236 5448 4264
rect 4571 4233 4583 4236
rect 4525 4227 4583 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 6086 4224 6092 4276
rect 6144 4224 6150 4276
rect 1857 4199 1915 4205
rect 1857 4165 1869 4199
rect 1903 4196 1915 4199
rect 1946 4196 1952 4208
rect 1903 4168 1952 4196
rect 1903 4165 1915 4168
rect 1857 4159 1915 4165
rect 1946 4156 1952 4168
rect 2004 4156 2010 4208
rect 3510 4196 3516 4208
rect 3082 4168 3516 4196
rect 3510 4156 3516 4168
rect 3568 4156 3574 4208
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 4120 4168 5488 4196
rect 4120 4156 4126 4168
rect 1578 4088 1584 4140
rect 1636 4088 1642 4140
rect 3694 4088 3700 4140
rect 3752 4088 3758 4140
rect 5460 4137 5488 4168
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4908 4100 4997 4128
rect 3786 4020 3792 4072
rect 3844 4020 3850 4072
rect 4246 4060 4252 4072
rect 3896 4032 4252 4060
rect 2866 3952 2872 4004
rect 2924 3992 2930 4004
rect 3896 3992 3924 4032
rect 4246 4020 4252 4032
rect 4304 4020 4310 4072
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 2924 3964 3924 3992
rect 4065 3995 4123 4001
rect 2924 3952 2930 3964
rect 4065 3961 4077 3995
rect 4111 3992 4123 3995
rect 4448 3992 4476 4023
rect 4908 4001 4936 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5491 4100 5733 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 5721 4097 5733 4100
rect 5767 4128 5779 4131
rect 6104 4128 6132 4224
rect 6454 4128 6460 4140
rect 5767 4100 6460 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4128 8815 4131
rect 10686 4128 10692 4140
rect 8803 4100 10692 4128
rect 8803 4097 8815 4100
rect 8757 4091 8815 4097
rect 10686 4088 10692 4100
rect 10744 4088 10750 4140
rect 4111 3964 4476 3992
rect 4893 3995 4951 4001
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 4893 3961 4905 3995
rect 4939 3961 4951 3995
rect 5534 3992 5540 4004
rect 4893 3955 4951 3961
rect 5184 3964 5540 3992
rect 3326 3884 3332 3936
rect 3384 3884 3390 3936
rect 5184 3933 5212 3964
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 5169 3927 5227 3933
rect 5169 3893 5181 3927
rect 5215 3893 5227 3927
rect 5169 3887 5227 3893
rect 5353 3927 5411 3933
rect 5353 3893 5365 3927
rect 5399 3924 5411 3927
rect 5442 3924 5448 3936
rect 5399 3896 5448 3924
rect 5399 3893 5411 3896
rect 5353 3887 5411 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3924 5687 3927
rect 6086 3924 6092 3936
rect 5675 3896 6092 3924
rect 5675 3893 5687 3896
rect 5629 3887 5687 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 8849 3927 8907 3933
rect 8849 3924 8861 3927
rect 8812 3896 8861 3924
rect 8812 3884 8818 3896
rect 8849 3893 8861 3896
rect 8895 3893 8907 3927
rect 8849 3887 8907 3893
rect 1104 3834 11868 3856
rect 1104 3782 2295 3834
rect 2347 3782 2359 3834
rect 2411 3782 2423 3834
rect 2475 3782 2487 3834
rect 2539 3782 2551 3834
rect 2603 3782 4986 3834
rect 5038 3782 5050 3834
rect 5102 3782 5114 3834
rect 5166 3782 5178 3834
rect 5230 3782 5242 3834
rect 5294 3782 7677 3834
rect 7729 3782 7741 3834
rect 7793 3782 7805 3834
rect 7857 3782 7869 3834
rect 7921 3782 7933 3834
rect 7985 3782 10368 3834
rect 10420 3782 10432 3834
rect 10484 3782 10496 3834
rect 10548 3782 10560 3834
rect 10612 3782 10624 3834
rect 10676 3782 11868 3834
rect 1104 3760 11868 3782
rect 3510 3680 3516 3732
rect 3568 3680 3574 3732
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 7650 3720 7656 3732
rect 7340 3692 7656 3720
rect 7340 3680 7346 3692
rect 7650 3680 7656 3692
rect 7708 3720 7714 3732
rect 7708 3692 9536 3720
rect 7708 3680 7714 3692
rect 2682 3652 2688 3664
rect 1780 3624 2688 3652
rect 1780 3525 1808 3624
rect 2682 3612 2688 3624
rect 2740 3612 2746 3664
rect 4893 3655 4951 3661
rect 4893 3621 4905 3655
rect 4939 3621 4951 3655
rect 4893 3615 4951 3621
rect 8941 3655 8999 3661
rect 8941 3621 8953 3655
rect 8987 3621 8999 3655
rect 8941 3615 8999 3621
rect 2038 3544 2044 3596
rect 2096 3544 2102 3596
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 4908 3584 4936 3615
rect 5994 3584 6000 3596
rect 4856 3556 6000 3584
rect 4856 3544 4862 3556
rect 5994 3544 6000 3556
rect 6052 3584 6058 3596
rect 6273 3587 6331 3593
rect 6273 3584 6285 3587
rect 6052 3556 6285 3584
rect 6052 3544 6058 3556
rect 6273 3553 6285 3556
rect 6319 3584 6331 3587
rect 7742 3584 7748 3596
rect 6319 3556 7748 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 7742 3544 7748 3556
rect 7800 3584 7806 3596
rect 7800 3556 8340 3584
rect 7800 3544 7806 3556
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 2130 3476 2136 3528
rect 2188 3516 2194 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 2188 3488 2237 3516
rect 2188 3476 2194 3488
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2961 3519 3019 3525
rect 2961 3516 2973 3519
rect 2225 3479 2283 3485
rect 2700 3488 2973 3516
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1397 3451 1455 3457
rect 1397 3448 1409 3451
rect 992 3420 1409 3448
rect 992 3408 998 3420
rect 1397 3417 1409 3420
rect 1443 3417 1455 3451
rect 1397 3411 1455 3417
rect 1854 3340 1860 3392
rect 1912 3380 1918 3392
rect 2314 3380 2320 3392
rect 1912 3352 2320 3380
rect 1912 3340 1918 3352
rect 2314 3340 2320 3352
rect 2372 3340 2378 3392
rect 2700 3389 2728 3488
rect 2961 3485 2973 3488
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 4062 3516 4068 3528
rect 3651 3488 4068 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 6178 3476 6184 3528
rect 6236 3476 6242 3528
rect 6546 3408 6552 3460
rect 6604 3408 6610 3460
rect 7282 3408 7288 3460
rect 7340 3408 7346 3460
rect 8202 3448 8208 3460
rect 8036 3420 8208 3448
rect 2685 3383 2743 3389
rect 2685 3349 2697 3383
rect 2731 3349 2743 3383
rect 2685 3343 2743 3349
rect 2774 3340 2780 3392
rect 2832 3340 2838 3392
rect 7834 3340 7840 3392
rect 7892 3380 7898 3392
rect 8036 3389 8064 3420
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 8312 3448 8340 3556
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 8956 3516 8984 3615
rect 9306 3612 9312 3664
rect 9364 3612 9370 3664
rect 9324 3584 9352 3612
rect 9508 3593 9536 3692
rect 8619 3488 8984 3516
rect 9048 3556 9352 3584
rect 9493 3587 9551 3593
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 9048 3448 9076 3556
rect 9493 3553 9505 3587
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 9582 3544 9588 3596
rect 9640 3544 9646 3596
rect 9122 3476 9128 3528
rect 9180 3516 9186 3528
rect 9306 3516 9312 3528
rect 9180 3488 9312 3516
rect 9180 3476 9186 3488
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3516 9459 3519
rect 9600 3516 9628 3544
rect 9447 3488 9628 3516
rect 9447 3485 9459 3488
rect 9401 3479 9459 3485
rect 8312 3420 9076 3448
rect 8021 3383 8079 3389
rect 8021 3380 8033 3383
rect 7892 3352 8033 3380
rect 7892 3340 7898 3352
rect 8021 3349 8033 3352
rect 8067 3349 8079 3383
rect 8021 3343 8079 3349
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8389 3383 8447 3389
rect 8389 3380 8401 3383
rect 8168 3352 8401 3380
rect 8168 3340 8174 3352
rect 8389 3349 8401 3352
rect 8435 3349 8447 3383
rect 8389 3343 8447 3349
rect 1104 3290 11868 3312
rect 1104 3238 2955 3290
rect 3007 3238 3019 3290
rect 3071 3238 3083 3290
rect 3135 3238 3147 3290
rect 3199 3238 3211 3290
rect 3263 3238 5646 3290
rect 5698 3238 5710 3290
rect 5762 3238 5774 3290
rect 5826 3238 5838 3290
rect 5890 3238 5902 3290
rect 5954 3238 8337 3290
rect 8389 3238 8401 3290
rect 8453 3238 8465 3290
rect 8517 3238 8529 3290
rect 8581 3238 8593 3290
rect 8645 3238 11028 3290
rect 11080 3238 11092 3290
rect 11144 3238 11156 3290
rect 11208 3238 11220 3290
rect 11272 3238 11284 3290
rect 11336 3238 11868 3290
rect 1104 3216 11868 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 4798 3176 4804 3188
rect 1636 3148 4804 3176
rect 1636 3136 1642 3148
rect 1688 3049 1716 3148
rect 3881 3111 3939 3117
rect 3881 3108 3893 3111
rect 3174 3080 3893 3108
rect 3881 3077 3893 3080
rect 3927 3077 3939 3111
rect 4062 3108 4068 3120
rect 3881 3071 3939 3077
rect 3996 3080 4068 3108
rect 3996 3049 4024 3080
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 4172 3049 4200 3148
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 6546 3136 6552 3188
rect 6604 3176 6610 3188
rect 6641 3179 6699 3185
rect 6641 3176 6653 3179
rect 6604 3148 6653 3176
rect 6604 3136 6610 3148
rect 6641 3145 6653 3148
rect 6687 3145 6699 3179
rect 6641 3139 6699 3145
rect 7377 3179 7435 3185
rect 7377 3145 7389 3179
rect 7423 3176 7435 3179
rect 7558 3176 7564 3188
rect 7423 3148 7564 3176
rect 7423 3145 7435 3148
rect 7377 3139 7435 3145
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 7834 3176 7840 3188
rect 7668 3148 7840 3176
rect 4433 3111 4491 3117
rect 4433 3077 4445 3111
rect 4479 3108 4491 3111
rect 4522 3108 4528 3120
rect 4479 3080 4528 3108
rect 4479 3077 4491 3080
rect 4433 3071 4491 3077
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 5442 3068 5448 3120
rect 5500 3068 5506 3120
rect 7190 3068 7196 3120
rect 7248 3108 7254 3120
rect 7285 3111 7343 3117
rect 7285 3108 7297 3111
rect 7248 3080 7297 3108
rect 7248 3068 7254 3080
rect 7285 3077 7297 3080
rect 7331 3108 7343 3111
rect 7668 3108 7696 3148
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9493 3179 9551 3185
rect 9493 3176 9505 3179
rect 9364 3148 9505 3176
rect 9364 3136 9370 3148
rect 9493 3145 9505 3148
rect 9539 3145 9551 3179
rect 9493 3139 9551 3145
rect 7331 3080 7696 3108
rect 7331 3077 7343 3080
rect 7285 3071 7343 3077
rect 8754 3068 8760 3120
rect 8812 3068 8818 3120
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3040 6883 3043
rect 7742 3040 7748 3052
rect 7800 3049 7806 3052
rect 6871 3012 6960 3040
rect 7710 3012 7748 3040
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2682 2972 2688 2984
rect 1995 2944 2688 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 3697 2975 3755 2981
rect 3697 2941 3709 2975
rect 3743 2972 3755 2975
rect 3743 2944 5856 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 2314 2796 2320 2848
rect 2372 2836 2378 2848
rect 3712 2836 3740 2935
rect 2372 2808 3740 2836
rect 5828 2836 5856 2944
rect 6178 2932 6184 2984
rect 6236 2932 6242 2984
rect 6932 2913 6960 3012
rect 7742 3000 7748 3012
rect 7800 3003 7810 3049
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 7800 3000 7806 3003
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 7650 2972 7656 2984
rect 7607 2944 7656 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8110 2972 8116 2984
rect 8067 2944 8116 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 6917 2907 6975 2913
rect 6917 2873 6929 2907
rect 6963 2873 6975 2907
rect 10980 2904 11008 3003
rect 6917 2867 6975 2873
rect 9048 2876 11008 2904
rect 9048 2836 9076 2876
rect 5828 2808 9076 2836
rect 2372 2796 2378 2808
rect 10686 2796 10692 2848
rect 10744 2836 10750 2848
rect 11057 2839 11115 2845
rect 11057 2836 11069 2839
rect 10744 2808 11069 2836
rect 10744 2796 10750 2808
rect 11057 2805 11069 2808
rect 11103 2805 11115 2839
rect 11057 2799 11115 2805
rect 1104 2746 11868 2768
rect 1104 2694 2295 2746
rect 2347 2694 2359 2746
rect 2411 2694 2423 2746
rect 2475 2694 2487 2746
rect 2539 2694 2551 2746
rect 2603 2694 4986 2746
rect 5038 2694 5050 2746
rect 5102 2694 5114 2746
rect 5166 2694 5178 2746
rect 5230 2694 5242 2746
rect 5294 2694 7677 2746
rect 7729 2694 7741 2746
rect 7793 2694 7805 2746
rect 7857 2694 7869 2746
rect 7921 2694 7933 2746
rect 7985 2694 10368 2746
rect 10420 2694 10432 2746
rect 10484 2694 10496 2746
rect 10548 2694 10560 2746
rect 10612 2694 10624 2746
rect 10676 2694 11868 2746
rect 1104 2672 11868 2694
rect 4540 2604 6224 2632
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2496 4031 2499
rect 4154 2496 4160 2508
rect 4019 2468 4160 2496
rect 4019 2465 4031 2468
rect 3973 2459 4031 2465
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 1854 2428 1860 2440
rect 1811 2400 1860 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 4540 2428 4568 2604
rect 6196 2576 6224 2604
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7340 2604 7389 2632
rect 7340 2592 7346 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 6178 2524 6184 2576
rect 6236 2524 6242 2576
rect 5718 2456 5724 2508
rect 5776 2456 5782 2508
rect 5994 2456 6000 2508
rect 6052 2456 6058 2508
rect 2915 2400 4568 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 6512 2400 7297 2428
rect 6512 2388 6518 2400
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 8202 2388 8208 2440
rect 8260 2428 8266 2440
rect 9033 2431 9091 2437
rect 9033 2428 9045 2431
rect 8260 2400 9045 2428
rect 8260 2388 8266 2400
rect 9033 2397 9045 2400
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 9490 2388 9496 2440
rect 9548 2388 9554 2440
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10836 2400 10977 2428
rect 10836 2388 10842 2400
rect 10965 2397 10977 2400
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 5290 2332 5396 2360
rect 1397 2323 1455 2329
rect 2590 2252 2596 2304
rect 2648 2252 2654 2304
rect 5368 2292 5396 2332
rect 5626 2320 5632 2372
rect 5684 2360 5690 2372
rect 6365 2363 6423 2369
rect 6365 2360 6377 2363
rect 5684 2332 6377 2360
rect 5684 2320 5690 2332
rect 6365 2329 6377 2332
rect 6411 2329 6423 2363
rect 6365 2323 6423 2329
rect 6733 2363 6791 2369
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 9508 2360 9536 2388
rect 6779 2332 9536 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 6086 2292 6092 2304
rect 5368 2264 6092 2292
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 8754 2252 8760 2304
rect 8812 2292 8818 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8812 2264 9137 2292
rect 8812 2252 8818 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 10870 2252 10876 2304
rect 10928 2292 10934 2304
rect 11057 2295 11115 2301
rect 11057 2292 11069 2295
rect 10928 2264 11069 2292
rect 10928 2252 10934 2264
rect 11057 2261 11069 2264
rect 11103 2261 11115 2295
rect 11057 2255 11115 2261
rect 1104 2202 11868 2224
rect 1104 2150 2955 2202
rect 3007 2150 3019 2202
rect 3071 2150 3083 2202
rect 3135 2150 3147 2202
rect 3199 2150 3211 2202
rect 3263 2150 5646 2202
rect 5698 2150 5710 2202
rect 5762 2150 5774 2202
rect 5826 2150 5838 2202
rect 5890 2150 5902 2202
rect 5954 2150 8337 2202
rect 8389 2150 8401 2202
rect 8453 2150 8465 2202
rect 8517 2150 8529 2202
rect 8581 2150 8593 2202
rect 8645 2150 11028 2202
rect 11080 2150 11092 2202
rect 11144 2150 11156 2202
rect 11208 2150 11220 2202
rect 11272 2150 11284 2202
rect 11336 2150 11868 2202
rect 1104 2128 11868 2150
rect 10686 1436 10692 1488
rect 10744 1476 10750 1488
rect 10962 1476 10968 1488
rect 10744 1448 10968 1476
rect 10744 1436 10750 1448
rect 10962 1436 10968 1448
rect 11020 1436 11026 1488
<< via1 >>
rect 2295 12486 2347 12538
rect 2359 12486 2411 12538
rect 2423 12486 2475 12538
rect 2487 12486 2539 12538
rect 2551 12486 2603 12538
rect 4986 12486 5038 12538
rect 5050 12486 5102 12538
rect 5114 12486 5166 12538
rect 5178 12486 5230 12538
rect 5242 12486 5294 12538
rect 7677 12486 7729 12538
rect 7741 12486 7793 12538
rect 7805 12486 7857 12538
rect 7869 12486 7921 12538
rect 7933 12486 7985 12538
rect 10368 12486 10420 12538
rect 10432 12486 10484 12538
rect 10496 12486 10548 12538
rect 10560 12486 10612 12538
rect 10624 12486 10676 12538
rect 1952 12384 2004 12436
rect 4712 12427 4764 12436
rect 4712 12393 4721 12427
rect 4721 12393 4755 12427
rect 4755 12393 4764 12427
rect 4712 12384 4764 12393
rect 10232 12384 10284 12436
rect 11244 12427 11296 12436
rect 11244 12393 11253 12427
rect 11253 12393 11287 12427
rect 11287 12393 11296 12427
rect 11244 12384 11296 12393
rect 8024 12359 8076 12368
rect 8024 12325 8033 12359
rect 8033 12325 8067 12359
rect 8067 12325 8076 12359
rect 8024 12316 8076 12325
rect 2228 12248 2280 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 1860 12180 1912 12232
rect 4712 12248 4764 12300
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 8668 12180 8720 12232
rect 11428 12180 11480 12232
rect 3424 12112 3476 12164
rect 4988 12155 5040 12164
rect 4988 12121 4997 12155
rect 4997 12121 5031 12155
rect 5031 12121 5040 12155
rect 4988 12112 5040 12121
rect 8116 12112 8168 12164
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 2780 12087 2832 12096
rect 2780 12053 2789 12087
rect 2789 12053 2823 12087
rect 2823 12053 2832 12087
rect 2780 12044 2832 12053
rect 8024 12044 8076 12096
rect 9036 12044 9088 12096
rect 2955 11942 3007 11994
rect 3019 11942 3071 11994
rect 3083 11942 3135 11994
rect 3147 11942 3199 11994
rect 3211 11942 3263 11994
rect 5646 11942 5698 11994
rect 5710 11942 5762 11994
rect 5774 11942 5826 11994
rect 5838 11942 5890 11994
rect 5902 11942 5954 11994
rect 8337 11942 8389 11994
rect 8401 11942 8453 11994
rect 8465 11942 8517 11994
rect 8529 11942 8581 11994
rect 8593 11942 8645 11994
rect 11028 11942 11080 11994
rect 11092 11942 11144 11994
rect 11156 11942 11208 11994
rect 11220 11942 11272 11994
rect 11284 11942 11336 11994
rect 2228 11840 2280 11892
rect 2780 11840 2832 11892
rect 940 11704 992 11756
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 2136 11500 2188 11509
rect 3700 11840 3752 11892
rect 4988 11840 5040 11892
rect 4068 11772 4120 11824
rect 6000 11772 6052 11824
rect 5356 11704 5408 11756
rect 8300 11704 8352 11756
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 4896 11636 4948 11688
rect 5540 11636 5592 11688
rect 9036 11840 9088 11892
rect 10140 11840 10192 11892
rect 9772 11772 9824 11824
rect 12900 11840 12952 11892
rect 2872 11500 2924 11552
rect 3240 11500 3292 11552
rect 3424 11500 3476 11552
rect 5448 11543 5500 11552
rect 5448 11509 5457 11543
rect 5457 11509 5491 11543
rect 5491 11509 5500 11543
rect 5448 11500 5500 11509
rect 5632 11500 5684 11552
rect 6644 11543 6696 11552
rect 6644 11509 6653 11543
rect 6653 11509 6687 11543
rect 6687 11509 6696 11543
rect 6644 11500 6696 11509
rect 8760 11500 8812 11552
rect 8852 11500 8904 11552
rect 9588 11500 9640 11552
rect 2295 11398 2347 11450
rect 2359 11398 2411 11450
rect 2423 11398 2475 11450
rect 2487 11398 2539 11450
rect 2551 11398 2603 11450
rect 4986 11398 5038 11450
rect 5050 11398 5102 11450
rect 5114 11398 5166 11450
rect 5178 11398 5230 11450
rect 5242 11398 5294 11450
rect 7677 11398 7729 11450
rect 7741 11398 7793 11450
rect 7805 11398 7857 11450
rect 7869 11398 7921 11450
rect 7933 11398 7985 11450
rect 10368 11398 10420 11450
rect 10432 11398 10484 11450
rect 10496 11398 10548 11450
rect 10560 11398 10612 11450
rect 10624 11398 10676 11450
rect 3240 11339 3292 11348
rect 3240 11305 3249 11339
rect 3249 11305 3283 11339
rect 3283 11305 3292 11339
rect 3240 11296 3292 11305
rect 4068 11296 4120 11348
rect 5632 11296 5684 11348
rect 8668 11296 8720 11348
rect 9772 11339 9824 11348
rect 9772 11305 9781 11339
rect 9781 11305 9815 11339
rect 9815 11305 9824 11339
rect 9772 11296 9824 11305
rect 2136 11160 2188 11212
rect 5540 11160 5592 11212
rect 8852 11160 8904 11212
rect 2412 11024 2464 11076
rect 3608 11092 3660 11144
rect 6644 11092 6696 11144
rect 8300 11092 8352 11144
rect 1860 10956 1912 11008
rect 2780 10956 2832 11008
rect 3332 10956 3384 11008
rect 3516 10956 3568 11008
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 7012 11067 7064 11076
rect 7012 11033 7021 11067
rect 7021 11033 7055 11067
rect 7055 11033 7064 11067
rect 7012 11024 7064 11033
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 9772 11024 9824 11076
rect 4712 10956 4764 11008
rect 5448 10956 5500 11008
rect 6000 10956 6052 11008
rect 6736 10956 6788 11008
rect 8760 10956 8812 11008
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 9956 10999 10008 11008
rect 9956 10965 9965 10999
rect 9965 10965 9999 10999
rect 9999 10965 10008 10999
rect 9956 10956 10008 10965
rect 2955 10854 3007 10906
rect 3019 10854 3071 10906
rect 3083 10854 3135 10906
rect 3147 10854 3199 10906
rect 3211 10854 3263 10906
rect 5646 10854 5698 10906
rect 5710 10854 5762 10906
rect 5774 10854 5826 10906
rect 5838 10854 5890 10906
rect 5902 10854 5954 10906
rect 8337 10854 8389 10906
rect 8401 10854 8453 10906
rect 8465 10854 8517 10906
rect 8529 10854 8581 10906
rect 8593 10854 8645 10906
rect 11028 10854 11080 10906
rect 11092 10854 11144 10906
rect 11156 10854 11208 10906
rect 11220 10854 11272 10906
rect 11284 10854 11336 10906
rect 2412 10795 2464 10804
rect 2412 10761 2421 10795
rect 2421 10761 2455 10795
rect 2455 10761 2464 10795
rect 2412 10752 2464 10761
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 3516 10752 3568 10804
rect 4528 10752 4580 10804
rect 5356 10752 5408 10804
rect 6000 10752 6052 10804
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 7012 10752 7064 10804
rect 11428 10752 11480 10804
rect 3056 10616 3108 10668
rect 3332 10659 3384 10668
rect 3332 10625 3341 10659
rect 3341 10625 3375 10659
rect 3375 10625 3384 10659
rect 3332 10616 3384 10625
rect 3516 10616 3568 10668
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 3700 10659 3752 10668
rect 3700 10625 3709 10659
rect 3709 10625 3743 10659
rect 3743 10625 3752 10659
rect 3700 10616 3752 10625
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 4712 10616 4764 10668
rect 4804 10659 4856 10668
rect 4804 10625 4813 10659
rect 4813 10625 4847 10659
rect 4847 10625 4856 10659
rect 4804 10616 4856 10625
rect 3148 10548 3200 10600
rect 4160 10548 4212 10600
rect 2780 10480 2832 10532
rect 3056 10523 3108 10532
rect 3056 10489 3065 10523
rect 3065 10489 3099 10523
rect 3099 10489 3108 10523
rect 3056 10480 3108 10489
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 5908 10548 5960 10557
rect 6828 10616 6880 10668
rect 4344 10480 4396 10532
rect 6644 10480 6696 10532
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 8944 10684 8996 10736
rect 9956 10684 10008 10736
rect 10876 10684 10928 10736
rect 7104 10548 7156 10600
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 8392 10659 8444 10668
rect 8392 10625 8401 10659
rect 8401 10625 8435 10659
rect 8435 10625 8444 10659
rect 8392 10616 8444 10625
rect 8668 10616 8720 10668
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 6736 10455 6788 10464
rect 6736 10421 6745 10455
rect 6745 10421 6779 10455
rect 6779 10421 6788 10455
rect 6736 10412 6788 10421
rect 8208 10480 8260 10532
rect 8300 10412 8352 10464
rect 9496 10412 9548 10464
rect 2295 10310 2347 10362
rect 2359 10310 2411 10362
rect 2423 10310 2475 10362
rect 2487 10310 2539 10362
rect 2551 10310 2603 10362
rect 4986 10310 5038 10362
rect 5050 10310 5102 10362
rect 5114 10310 5166 10362
rect 5178 10310 5230 10362
rect 5242 10310 5294 10362
rect 7677 10310 7729 10362
rect 7741 10310 7793 10362
rect 7805 10310 7857 10362
rect 7869 10310 7921 10362
rect 7933 10310 7985 10362
rect 10368 10310 10420 10362
rect 10432 10310 10484 10362
rect 10496 10310 10548 10362
rect 10560 10310 10612 10362
rect 10624 10310 10676 10362
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 3608 10208 3660 10260
rect 3700 10208 3752 10260
rect 3976 10208 4028 10260
rect 4528 10208 4580 10260
rect 3056 10140 3108 10192
rect 3516 10140 3568 10192
rect 5908 10251 5960 10260
rect 5908 10217 5917 10251
rect 5917 10217 5951 10251
rect 5951 10217 5960 10251
rect 5908 10208 5960 10217
rect 6828 10208 6880 10260
rect 7380 10208 7432 10260
rect 10140 10208 10192 10260
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 7104 10140 7156 10192
rect 1860 10004 1912 10056
rect 2504 10004 2556 10056
rect 3884 10072 3936 10124
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 6736 10072 6788 10124
rect 2688 9936 2740 9988
rect 4068 10004 4120 10056
rect 3700 9936 3752 9988
rect 4804 10004 4856 10056
rect 8392 10140 8444 10192
rect 9312 10140 9364 10192
rect 1584 9868 1636 9920
rect 4252 9868 4304 9920
rect 4896 9868 4948 9920
rect 6920 9868 6972 9920
rect 8208 10072 8260 10124
rect 8760 10072 8812 10124
rect 9864 10140 9916 10192
rect 9772 10072 9824 10124
rect 8300 10004 8352 10056
rect 10692 10004 10744 10056
rect 9956 9936 10008 9988
rect 11428 10004 11480 10056
rect 11520 9936 11572 9988
rect 8668 9868 8720 9920
rect 9680 9868 9732 9920
rect 2955 9766 3007 9818
rect 3019 9766 3071 9818
rect 3083 9766 3135 9818
rect 3147 9766 3199 9818
rect 3211 9766 3263 9818
rect 5646 9766 5698 9818
rect 5710 9766 5762 9818
rect 5774 9766 5826 9818
rect 5838 9766 5890 9818
rect 5902 9766 5954 9818
rect 8337 9766 8389 9818
rect 8401 9766 8453 9818
rect 8465 9766 8517 9818
rect 8529 9766 8581 9818
rect 8593 9766 8645 9818
rect 11028 9766 11080 9818
rect 11092 9766 11144 9818
rect 11156 9766 11208 9818
rect 11220 9766 11272 9818
rect 11284 9766 11336 9818
rect 2688 9596 2740 9648
rect 5540 9596 5592 9648
rect 7012 9596 7064 9648
rect 9128 9596 9180 9648
rect 9772 9664 9824 9716
rect 9956 9664 10008 9716
rect 12072 9664 12124 9716
rect 9312 9639 9364 9648
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 3424 9528 3476 9580
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 8944 9460 8996 9469
rect 9680 9460 9732 9512
rect 8852 9392 8904 9444
rect 3608 9324 3660 9376
rect 8760 9324 8812 9376
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 9956 9324 10008 9376
rect 11520 9324 11572 9376
rect 2295 9222 2347 9274
rect 2359 9222 2411 9274
rect 2423 9222 2475 9274
rect 2487 9222 2539 9274
rect 2551 9222 2603 9274
rect 4986 9222 5038 9274
rect 5050 9222 5102 9274
rect 5114 9222 5166 9274
rect 5178 9222 5230 9274
rect 5242 9222 5294 9274
rect 7677 9222 7729 9274
rect 7741 9222 7793 9274
rect 7805 9222 7857 9274
rect 7869 9222 7921 9274
rect 7933 9222 7985 9274
rect 10368 9222 10420 9274
rect 10432 9222 10484 9274
rect 10496 9222 10548 9274
rect 10560 9222 10612 9274
rect 10624 9222 10676 9274
rect 4160 9120 4212 9172
rect 4712 9120 4764 9172
rect 5356 9120 5408 9172
rect 8852 9120 8904 9172
rect 9680 9120 9732 9172
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 940 8916 992 8968
rect 2044 8891 2096 8900
rect 2044 8857 2053 8891
rect 2053 8857 2087 8891
rect 2087 8857 2096 8891
rect 2044 8848 2096 8857
rect 3516 8916 3568 8968
rect 3700 8916 3752 8968
rect 3884 8916 3936 8968
rect 8944 9052 8996 9104
rect 9404 9052 9456 9104
rect 9496 9052 9548 9104
rect 6368 8984 6420 9036
rect 7012 8984 7064 9036
rect 8760 9027 8812 9036
rect 8760 8993 8769 9027
rect 8769 8993 8803 9027
rect 8803 8993 8812 9027
rect 8760 8984 8812 8993
rect 2780 8780 2832 8832
rect 2872 8823 2924 8832
rect 2872 8789 2881 8823
rect 2881 8789 2915 8823
rect 2915 8789 2924 8823
rect 2872 8780 2924 8789
rect 3332 8780 3384 8832
rect 4528 8891 4580 8900
rect 4528 8857 4537 8891
rect 4537 8857 4571 8891
rect 4571 8857 4580 8891
rect 4528 8848 4580 8857
rect 4620 8891 4672 8900
rect 4620 8857 4629 8891
rect 4629 8857 4663 8891
rect 4663 8857 4672 8891
rect 4620 8848 4672 8857
rect 5172 8891 5224 8900
rect 5172 8857 5181 8891
rect 5181 8857 5215 8891
rect 5215 8857 5224 8891
rect 5172 8848 5224 8857
rect 6184 8848 6236 8900
rect 8852 8916 8904 8968
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 9772 8984 9824 9036
rect 7104 8780 7156 8832
rect 8944 8780 8996 8832
rect 10140 8848 10192 8900
rect 9956 8780 10008 8832
rect 2955 8678 3007 8730
rect 3019 8678 3071 8730
rect 3083 8678 3135 8730
rect 3147 8678 3199 8730
rect 3211 8678 3263 8730
rect 5646 8678 5698 8730
rect 5710 8678 5762 8730
rect 5774 8678 5826 8730
rect 5838 8678 5890 8730
rect 5902 8678 5954 8730
rect 8337 8678 8389 8730
rect 8401 8678 8453 8730
rect 8465 8678 8517 8730
rect 8529 8678 8581 8730
rect 8593 8678 8645 8730
rect 11028 8678 11080 8730
rect 11092 8678 11144 8730
rect 11156 8678 11208 8730
rect 11220 8678 11272 8730
rect 11284 8678 11336 8730
rect 2872 8576 2924 8628
rect 3332 8576 3384 8628
rect 4620 8576 4672 8628
rect 4712 8619 4764 8628
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 6184 8576 6236 8628
rect 1768 8440 1820 8492
rect 3424 8508 3476 8560
rect 2964 8372 3016 8424
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 6552 8508 6604 8560
rect 7104 8508 7156 8560
rect 8852 8508 8904 8560
rect 8944 8508 8996 8560
rect 2228 8304 2280 8356
rect 3700 8304 3752 8356
rect 4252 8372 4304 8424
rect 4620 8415 4672 8424
rect 4620 8381 4629 8415
rect 4629 8381 4663 8415
rect 4663 8381 4672 8415
rect 4620 8372 4672 8381
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 6092 8372 6144 8424
rect 7012 8372 7064 8424
rect 8024 8304 8076 8356
rect 10140 8576 10192 8628
rect 10784 8576 10836 8628
rect 10876 8508 10928 8560
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9588 8483 9640 8492
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 9588 8440 9640 8449
rect 10232 8372 10284 8424
rect 3792 8236 3844 8288
rect 9864 8236 9916 8288
rect 2295 8134 2347 8186
rect 2359 8134 2411 8186
rect 2423 8134 2475 8186
rect 2487 8134 2539 8186
rect 2551 8134 2603 8186
rect 4986 8134 5038 8186
rect 5050 8134 5102 8186
rect 5114 8134 5166 8186
rect 5178 8134 5230 8186
rect 5242 8134 5294 8186
rect 7677 8134 7729 8186
rect 7741 8134 7793 8186
rect 7805 8134 7857 8186
rect 7869 8134 7921 8186
rect 7933 8134 7985 8186
rect 10368 8134 10420 8186
rect 10432 8134 10484 8186
rect 10496 8134 10548 8186
rect 10560 8134 10612 8186
rect 10624 8134 10676 8186
rect 6368 8032 6420 8084
rect 9036 8032 9088 8084
rect 9680 8032 9732 8084
rect 9956 8032 10008 8084
rect 10232 8032 10284 8084
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 1952 7896 2004 7948
rect 3516 7896 3568 7948
rect 8024 7896 8076 7948
rect 2044 7828 2096 7880
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 8668 7896 8720 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 9864 7939 9916 7948
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 9128 7828 9180 7880
rect 1768 7803 1820 7812
rect 1768 7769 1777 7803
rect 1777 7769 1811 7803
rect 1811 7769 1820 7803
rect 1768 7760 1820 7769
rect 6920 7760 6972 7812
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 7288 7692 7340 7744
rect 10692 7964 10744 8016
rect 10784 7692 10836 7744
rect 2955 7590 3007 7642
rect 3019 7590 3071 7642
rect 3083 7590 3135 7642
rect 3147 7590 3199 7642
rect 3211 7590 3263 7642
rect 5646 7590 5698 7642
rect 5710 7590 5762 7642
rect 5774 7590 5826 7642
rect 5838 7590 5890 7642
rect 5902 7590 5954 7642
rect 8337 7590 8389 7642
rect 8401 7590 8453 7642
rect 8465 7590 8517 7642
rect 8529 7590 8581 7642
rect 8593 7590 8645 7642
rect 11028 7590 11080 7642
rect 11092 7590 11144 7642
rect 11156 7590 11208 7642
rect 11220 7590 11272 7642
rect 11284 7590 11336 7642
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 3424 7488 3476 7540
rect 3792 7420 3844 7472
rect 3516 7352 3568 7404
rect 8208 7352 8260 7404
rect 3332 7284 3384 7336
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 3884 7284 3936 7336
rect 4620 7284 4672 7336
rect 4160 7148 4212 7200
rect 5540 7148 5592 7200
rect 6920 7148 6972 7200
rect 2295 7046 2347 7098
rect 2359 7046 2411 7098
rect 2423 7046 2475 7098
rect 2487 7046 2539 7098
rect 2551 7046 2603 7098
rect 4986 7046 5038 7098
rect 5050 7046 5102 7098
rect 5114 7046 5166 7098
rect 5178 7046 5230 7098
rect 5242 7046 5294 7098
rect 7677 7046 7729 7098
rect 7741 7046 7793 7098
rect 7805 7046 7857 7098
rect 7869 7046 7921 7098
rect 7933 7046 7985 7098
rect 10368 7046 10420 7098
rect 10432 7046 10484 7098
rect 10496 7046 10548 7098
rect 10560 7046 10612 7098
rect 10624 7046 10676 7098
rect 3608 6987 3660 6996
rect 3608 6953 3617 6987
rect 3617 6953 3651 6987
rect 3651 6953 3660 6987
rect 3608 6944 3660 6953
rect 6828 6944 6880 6996
rect 3424 6876 3476 6928
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 2044 6808 2096 6860
rect 1676 6740 1728 6792
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 3516 6740 3568 6792
rect 2228 6604 2280 6656
rect 3332 6604 3384 6656
rect 5356 6740 5408 6792
rect 3884 6672 3936 6724
rect 5172 6672 5224 6724
rect 9680 6876 9732 6928
rect 6828 6740 6880 6792
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 7288 6740 7340 6792
rect 7380 6740 7432 6792
rect 9588 6808 9640 6860
rect 7472 6715 7524 6724
rect 7472 6681 7481 6715
rect 7481 6681 7515 6715
rect 7515 6681 7524 6715
rect 7472 6672 7524 6681
rect 8760 6740 8812 6792
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9220 6740 9272 6792
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 9496 6672 9548 6724
rect 6000 6604 6052 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 6552 6604 6604 6656
rect 7288 6647 7340 6656
rect 7288 6613 7315 6647
rect 7315 6613 7340 6647
rect 7288 6604 7340 6613
rect 7564 6604 7616 6656
rect 8852 6604 8904 6656
rect 9404 6604 9456 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 2955 6502 3007 6554
rect 3019 6502 3071 6554
rect 3083 6502 3135 6554
rect 3147 6502 3199 6554
rect 3211 6502 3263 6554
rect 5646 6502 5698 6554
rect 5710 6502 5762 6554
rect 5774 6502 5826 6554
rect 5838 6502 5890 6554
rect 5902 6502 5954 6554
rect 8337 6502 8389 6554
rect 8401 6502 8453 6554
rect 8465 6502 8517 6554
rect 8529 6502 8581 6554
rect 8593 6502 8645 6554
rect 11028 6502 11080 6554
rect 11092 6502 11144 6554
rect 11156 6502 11208 6554
rect 11220 6502 11272 6554
rect 11284 6502 11336 6554
rect 2228 6400 2280 6452
rect 3516 6400 3568 6452
rect 3884 6443 3936 6452
rect 3884 6409 3893 6443
rect 3893 6409 3927 6443
rect 3927 6409 3936 6443
rect 3884 6400 3936 6409
rect 4528 6400 4580 6452
rect 2044 6264 2096 6316
rect 4436 6332 4488 6384
rect 5080 6400 5132 6452
rect 5172 6443 5224 6452
rect 5172 6409 5181 6443
rect 5181 6409 5215 6443
rect 5215 6409 5224 6443
rect 5172 6400 5224 6409
rect 6000 6400 6052 6452
rect 7012 6400 7064 6452
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 6276 6332 6328 6384
rect 4344 6264 4396 6273
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 5356 6264 5408 6316
rect 5540 6264 5592 6316
rect 2688 6128 2740 6180
rect 2964 6171 3016 6180
rect 2964 6137 2973 6171
rect 2973 6137 3007 6171
rect 3007 6137 3016 6171
rect 2964 6128 3016 6137
rect 5080 6128 5132 6180
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 8944 6400 8996 6452
rect 9496 6400 9548 6452
rect 9680 6400 9732 6452
rect 6828 6196 6880 6248
rect 7104 6196 7156 6248
rect 8024 6264 8076 6316
rect 8484 6332 8536 6384
rect 8300 6264 8352 6316
rect 9312 6264 9364 6316
rect 10876 6264 10928 6316
rect 8208 6196 8260 6248
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 9036 6239 9088 6248
rect 9036 6205 9045 6239
rect 9045 6205 9079 6239
rect 9079 6205 9088 6239
rect 9036 6196 9088 6205
rect 9496 6239 9548 6248
rect 9496 6205 9505 6239
rect 9505 6205 9539 6239
rect 9539 6205 9548 6239
rect 9496 6196 9548 6205
rect 9772 6196 9824 6248
rect 4436 6103 4488 6112
rect 4436 6069 4445 6103
rect 4445 6069 4479 6103
rect 4479 6069 4488 6103
rect 4436 6060 4488 6069
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 5540 6103 5592 6112
rect 5540 6069 5549 6103
rect 5549 6069 5583 6103
rect 5583 6069 5592 6103
rect 5540 6060 5592 6069
rect 5632 6103 5684 6112
rect 5632 6069 5641 6103
rect 5641 6069 5675 6103
rect 5675 6069 5684 6103
rect 5632 6060 5684 6069
rect 7012 6060 7064 6112
rect 8484 6060 8536 6112
rect 9036 6060 9088 6112
rect 9312 6060 9364 6112
rect 2295 5958 2347 6010
rect 2359 5958 2411 6010
rect 2423 5958 2475 6010
rect 2487 5958 2539 6010
rect 2551 5958 2603 6010
rect 4986 5958 5038 6010
rect 5050 5958 5102 6010
rect 5114 5958 5166 6010
rect 5178 5958 5230 6010
rect 5242 5958 5294 6010
rect 7677 5958 7729 6010
rect 7741 5958 7793 6010
rect 7805 5958 7857 6010
rect 7869 5958 7921 6010
rect 7933 5958 7985 6010
rect 10368 5958 10420 6010
rect 10432 5958 10484 6010
rect 10496 5958 10548 6010
rect 10560 5958 10612 6010
rect 10624 5958 10676 6010
rect 1860 5856 1912 5908
rect 3884 5856 3936 5908
rect 4344 5856 4396 5908
rect 4712 5856 4764 5908
rect 5080 5856 5132 5908
rect 6920 5856 6972 5908
rect 8116 5856 8168 5908
rect 8668 5856 8720 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 9220 5856 9272 5908
rect 9864 5856 9916 5908
rect 10692 5856 10744 5908
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 3332 5720 3384 5772
rect 2596 5652 2648 5704
rect 4160 5763 4212 5772
rect 4160 5729 4169 5763
rect 4169 5729 4203 5763
rect 4203 5729 4212 5763
rect 4160 5720 4212 5729
rect 4896 5720 4948 5772
rect 6828 5788 6880 5840
rect 5632 5720 5684 5772
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 6276 5652 6328 5704
rect 8576 5720 8628 5772
rect 8116 5652 8168 5704
rect 8208 5652 8260 5704
rect 8852 5720 8904 5772
rect 9036 5763 9088 5772
rect 9036 5729 9045 5763
rect 9045 5729 9079 5763
rect 9079 5729 9088 5763
rect 9036 5720 9088 5729
rect 9312 5720 9364 5772
rect 9588 5720 9640 5772
rect 2964 5516 3016 5568
rect 3700 5516 3752 5568
rect 4528 5559 4580 5568
rect 4528 5525 4537 5559
rect 4537 5525 4571 5559
rect 4571 5525 4580 5559
rect 4528 5516 4580 5525
rect 7104 5584 7156 5636
rect 9496 5652 9548 5704
rect 8852 5584 8904 5636
rect 9772 5584 9824 5636
rect 11796 5652 11848 5704
rect 5540 5516 5592 5568
rect 8944 5516 8996 5568
rect 9404 5516 9456 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 2955 5414 3007 5466
rect 3019 5414 3071 5466
rect 3083 5414 3135 5466
rect 3147 5414 3199 5466
rect 3211 5414 3263 5466
rect 5646 5414 5698 5466
rect 5710 5414 5762 5466
rect 5774 5414 5826 5466
rect 5838 5414 5890 5466
rect 5902 5414 5954 5466
rect 8337 5414 8389 5466
rect 8401 5414 8453 5466
rect 8465 5414 8517 5466
rect 8529 5414 8581 5466
rect 8593 5414 8645 5466
rect 11028 5414 11080 5466
rect 11092 5414 11144 5466
rect 11156 5414 11208 5466
rect 11220 5414 11272 5466
rect 11284 5414 11336 5466
rect 2688 5312 2740 5364
rect 4712 5355 4764 5364
rect 4712 5321 4721 5355
rect 4721 5321 4755 5355
rect 4755 5321 4764 5355
rect 4712 5312 4764 5321
rect 4896 5312 4948 5364
rect 9128 5312 9180 5364
rect 9404 5312 9456 5364
rect 940 5244 992 5296
rect 1676 5244 1728 5296
rect 3332 5244 3384 5296
rect 2044 5108 2096 5160
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 4436 5108 4488 5160
rect 9036 5244 9088 5296
rect 5356 5176 5408 5228
rect 6828 5176 6880 5228
rect 7288 5176 7340 5228
rect 8760 5176 8812 5228
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 9588 5083 9640 5092
rect 9588 5049 9597 5083
rect 9597 5049 9631 5083
rect 9631 5049 9640 5083
rect 9588 5040 9640 5049
rect 2872 4972 2924 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 2295 4870 2347 4922
rect 2359 4870 2411 4922
rect 2423 4870 2475 4922
rect 2487 4870 2539 4922
rect 2551 4870 2603 4922
rect 4986 4870 5038 4922
rect 5050 4870 5102 4922
rect 5114 4870 5166 4922
rect 5178 4870 5230 4922
rect 5242 4870 5294 4922
rect 7677 4870 7729 4922
rect 7741 4870 7793 4922
rect 7805 4870 7857 4922
rect 7869 4870 7921 4922
rect 7933 4870 7985 4922
rect 10368 4870 10420 4922
rect 10432 4870 10484 4922
rect 10496 4870 10548 4922
rect 10560 4870 10612 4922
rect 10624 4870 10676 4922
rect 1952 4768 2004 4820
rect 5540 4768 5592 4820
rect 9220 4768 9272 4820
rect 7104 4700 7156 4752
rect 4436 4675 4488 4684
rect 4436 4641 4445 4675
rect 4445 4641 4479 4675
rect 4479 4641 4488 4675
rect 4436 4632 4488 4641
rect 6828 4632 6880 4684
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 8760 4700 8812 4752
rect 8852 4632 8904 4684
rect 8668 4564 8720 4616
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 1952 4471 2004 4480
rect 1952 4437 1961 4471
rect 1961 4437 1995 4471
rect 1995 4437 2004 4471
rect 1952 4428 2004 4437
rect 3792 4428 3844 4480
rect 7196 4428 7248 4480
rect 7564 4471 7616 4480
rect 7564 4437 7573 4471
rect 7573 4437 7607 4471
rect 7607 4437 7616 4471
rect 7564 4428 7616 4437
rect 9588 4471 9640 4480
rect 9588 4437 9597 4471
rect 9597 4437 9631 4471
rect 9631 4437 9640 4471
rect 9588 4428 9640 4437
rect 2955 4326 3007 4378
rect 3019 4326 3071 4378
rect 3083 4326 3135 4378
rect 3147 4326 3199 4378
rect 3211 4326 3263 4378
rect 5646 4326 5698 4378
rect 5710 4326 5762 4378
rect 5774 4326 5826 4378
rect 5838 4326 5890 4378
rect 5902 4326 5954 4378
rect 8337 4326 8389 4378
rect 8401 4326 8453 4378
rect 8465 4326 8517 4378
rect 8529 4326 8581 4378
rect 8593 4326 8645 4378
rect 11028 4326 11080 4378
rect 11092 4326 11144 4378
rect 11156 4326 11208 4378
rect 11220 4326 11272 4378
rect 11284 4326 11336 4378
rect 2688 4224 2740 4276
rect 4160 4224 4212 4276
rect 5448 4224 5500 4276
rect 6092 4224 6144 4276
rect 1952 4156 2004 4208
rect 3516 4156 3568 4208
rect 4068 4156 4120 4208
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 4252 4063 4304 4072
rect 2872 3952 2924 4004
rect 4252 4029 4261 4063
rect 4261 4029 4295 4063
rect 4295 4029 4304 4063
rect 4252 4020 4304 4029
rect 6460 4088 6512 4140
rect 10692 4088 10744 4140
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 3332 3884 3384 3893
rect 5540 3952 5592 4004
rect 5448 3884 5500 3936
rect 6092 3884 6144 3936
rect 8760 3884 8812 3936
rect 2295 3782 2347 3834
rect 2359 3782 2411 3834
rect 2423 3782 2475 3834
rect 2487 3782 2539 3834
rect 2551 3782 2603 3834
rect 4986 3782 5038 3834
rect 5050 3782 5102 3834
rect 5114 3782 5166 3834
rect 5178 3782 5230 3834
rect 5242 3782 5294 3834
rect 7677 3782 7729 3834
rect 7741 3782 7793 3834
rect 7805 3782 7857 3834
rect 7869 3782 7921 3834
rect 7933 3782 7985 3834
rect 10368 3782 10420 3834
rect 10432 3782 10484 3834
rect 10496 3782 10548 3834
rect 10560 3782 10612 3834
rect 10624 3782 10676 3834
rect 3516 3723 3568 3732
rect 3516 3689 3525 3723
rect 3525 3689 3559 3723
rect 3559 3689 3568 3723
rect 3516 3680 3568 3689
rect 7288 3680 7340 3732
rect 7656 3680 7708 3732
rect 2688 3612 2740 3664
rect 2044 3587 2096 3596
rect 2044 3553 2053 3587
rect 2053 3553 2087 3587
rect 2087 3553 2096 3587
rect 2044 3544 2096 3553
rect 4804 3544 4856 3596
rect 6000 3544 6052 3596
rect 7748 3544 7800 3596
rect 2136 3476 2188 3528
rect 940 3408 992 3460
rect 1860 3340 1912 3392
rect 2320 3383 2372 3392
rect 2320 3349 2329 3383
rect 2329 3349 2363 3383
rect 2363 3349 2372 3383
rect 2320 3340 2372 3349
rect 4068 3476 4120 3528
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 6552 3451 6604 3460
rect 6552 3417 6561 3451
rect 6561 3417 6595 3451
rect 6595 3417 6604 3451
rect 6552 3408 6604 3417
rect 7288 3408 7340 3460
rect 2780 3383 2832 3392
rect 2780 3349 2789 3383
rect 2789 3349 2823 3383
rect 2823 3349 2832 3383
rect 2780 3340 2832 3349
rect 7840 3340 7892 3392
rect 8208 3408 8260 3460
rect 9312 3612 9364 3664
rect 9588 3544 9640 3596
rect 9128 3476 9180 3528
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 8116 3340 8168 3392
rect 2955 3238 3007 3290
rect 3019 3238 3071 3290
rect 3083 3238 3135 3290
rect 3147 3238 3199 3290
rect 3211 3238 3263 3290
rect 5646 3238 5698 3290
rect 5710 3238 5762 3290
rect 5774 3238 5826 3290
rect 5838 3238 5890 3290
rect 5902 3238 5954 3290
rect 8337 3238 8389 3290
rect 8401 3238 8453 3290
rect 8465 3238 8517 3290
rect 8529 3238 8581 3290
rect 8593 3238 8645 3290
rect 11028 3238 11080 3290
rect 11092 3238 11144 3290
rect 11156 3238 11208 3290
rect 11220 3238 11272 3290
rect 11284 3238 11336 3290
rect 1584 3136 1636 3188
rect 4068 3068 4120 3120
rect 4804 3136 4856 3188
rect 6552 3136 6604 3188
rect 7564 3136 7616 3188
rect 4528 3068 4580 3120
rect 5448 3068 5500 3120
rect 7196 3068 7248 3120
rect 7840 3136 7892 3188
rect 9312 3136 9364 3188
rect 8760 3068 8812 3120
rect 7748 3043 7800 3052
rect 2688 2932 2740 2984
rect 2320 2796 2372 2848
rect 6184 2975 6236 2984
rect 6184 2941 6193 2975
rect 6193 2941 6227 2975
rect 6227 2941 6236 2975
rect 6184 2932 6236 2941
rect 7748 3009 7764 3043
rect 7764 3009 7798 3043
rect 7798 3009 7800 3043
rect 7748 3000 7800 3009
rect 7656 2932 7708 2984
rect 8116 2932 8168 2984
rect 10692 2796 10744 2848
rect 2295 2694 2347 2746
rect 2359 2694 2411 2746
rect 2423 2694 2475 2746
rect 2487 2694 2539 2746
rect 2551 2694 2603 2746
rect 4986 2694 5038 2746
rect 5050 2694 5102 2746
rect 5114 2694 5166 2746
rect 5178 2694 5230 2746
rect 5242 2694 5294 2746
rect 7677 2694 7729 2746
rect 7741 2694 7793 2746
rect 7805 2694 7857 2746
rect 7869 2694 7921 2746
rect 7933 2694 7985 2746
rect 10368 2694 10420 2746
rect 10432 2694 10484 2746
rect 10496 2694 10548 2746
rect 10560 2694 10612 2746
rect 10624 2694 10676 2746
rect 4160 2456 4212 2508
rect 1860 2388 1912 2440
rect 7288 2592 7340 2644
rect 6184 2524 6236 2576
rect 5724 2499 5776 2508
rect 5724 2465 5733 2499
rect 5733 2465 5767 2499
rect 5767 2465 5776 2499
rect 5724 2456 5776 2465
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 6460 2388 6512 2440
rect 8208 2388 8260 2440
rect 9496 2388 9548 2440
rect 10784 2388 10836 2440
rect 20 2320 72 2372
rect 2596 2295 2648 2304
rect 2596 2261 2605 2295
rect 2605 2261 2639 2295
rect 2639 2261 2648 2295
rect 2596 2252 2648 2261
rect 5632 2320 5684 2372
rect 6092 2252 6144 2304
rect 8760 2252 8812 2304
rect 10876 2252 10928 2304
rect 2955 2150 3007 2202
rect 3019 2150 3071 2202
rect 3083 2150 3135 2202
rect 3147 2150 3199 2202
rect 3211 2150 3263 2202
rect 5646 2150 5698 2202
rect 5710 2150 5762 2202
rect 5774 2150 5826 2202
rect 5838 2150 5890 2202
rect 5902 2150 5954 2202
rect 8337 2150 8389 2202
rect 8401 2150 8453 2202
rect 8465 2150 8517 2202
rect 8529 2150 8581 2202
rect 8593 2150 8645 2202
rect 11028 2150 11080 2202
rect 11092 2150 11144 2202
rect 11156 2150 11208 2202
rect 11220 2150 11272 2202
rect 11284 2150 11336 2202
rect 10692 1436 10744 1488
rect 10968 1436 11020 1488
<< metal2 >>
rect 1950 14346 2006 15146
rect 4526 14346 4582 15146
rect 7746 14498 7802 15146
rect 10322 14498 10378 15146
rect 7746 14470 8064 14498
rect 7746 14346 7802 14470
rect 1398 14104 1454 14113
rect 1398 14039 1454 14048
rect 1412 12238 1440 14039
rect 1964 12442 1992 14346
rect 2295 12540 2603 12549
rect 2295 12538 2301 12540
rect 2357 12538 2381 12540
rect 2437 12538 2461 12540
rect 2517 12538 2541 12540
rect 2597 12538 2603 12540
rect 2357 12486 2359 12538
rect 2539 12486 2541 12538
rect 2295 12484 2301 12486
rect 2357 12484 2381 12486
rect 2437 12484 2461 12486
rect 2517 12484 2541 12486
rect 2597 12484 2603 12486
rect 2295 12475 2603 12484
rect 1952 12436 2004 12442
rect 4540 12434 4568 14346
rect 4986 12540 5294 12549
rect 4986 12538 4992 12540
rect 5048 12538 5072 12540
rect 5128 12538 5152 12540
rect 5208 12538 5232 12540
rect 5288 12538 5294 12540
rect 5048 12486 5050 12538
rect 5230 12486 5232 12538
rect 4986 12484 4992 12486
rect 5048 12484 5072 12486
rect 5128 12484 5152 12486
rect 5208 12484 5232 12486
rect 5288 12484 5294 12486
rect 4986 12475 5294 12484
rect 7677 12540 7985 12549
rect 7677 12538 7683 12540
rect 7739 12538 7763 12540
rect 7819 12538 7843 12540
rect 7899 12538 7923 12540
rect 7979 12538 7985 12540
rect 7739 12486 7741 12538
rect 7921 12486 7923 12538
rect 7677 12484 7683 12486
rect 7739 12484 7763 12486
rect 7819 12484 7843 12486
rect 7899 12484 7923 12486
rect 7979 12484 7985 12486
rect 7677 12475 7985 12484
rect 4712 12436 4764 12442
rect 4540 12406 4712 12434
rect 1952 12378 2004 12384
rect 4712 12378 4764 12384
rect 8036 12374 8064 14470
rect 10244 14470 10378 14498
rect 10244 12442 10272 14470
rect 10322 14346 10378 14470
rect 12898 14346 12954 15146
rect 10368 12540 10676 12549
rect 10368 12538 10374 12540
rect 10430 12538 10454 12540
rect 10510 12538 10534 12540
rect 10590 12538 10614 12540
rect 10670 12538 10676 12540
rect 10430 12486 10432 12538
rect 10612 12486 10614 12538
rect 10368 12484 10374 12486
rect 10430 12484 10454 12486
rect 10510 12484 10534 12486
rect 10590 12484 10614 12486
rect 10670 12484 10676 12486
rect 10368 12475 10676 12484
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 8024 12368 8076 12374
rect 11256 12345 11284 12378
rect 8024 12310 8076 12316
rect 11242 12336 11298 12345
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 10140 12300 10192 12306
rect 11242 12271 11298 12280
rect 10140 12242 10192 12248
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 1596 9926 1624 12038
rect 1872 11014 1900 12174
rect 2240 11898 2268 12242
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2792 11898 2820 12038
rect 2955 11996 3263 12005
rect 2955 11994 2961 11996
rect 3017 11994 3041 11996
rect 3097 11994 3121 11996
rect 3177 11994 3201 11996
rect 3257 11994 3263 11996
rect 3017 11942 3019 11994
rect 3199 11942 3201 11994
rect 2955 11940 2961 11942
rect 3017 11940 3041 11942
rect 3097 11940 3121 11942
rect 3177 11940 3201 11942
rect 3257 11940 3263 11942
rect 2955 11931 3263 11940
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 3436 11558 3464 12106
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 2148 11218 2176 11494
rect 2295 11452 2603 11461
rect 2295 11450 2301 11452
rect 2357 11450 2381 11452
rect 2437 11450 2461 11452
rect 2517 11450 2541 11452
rect 2597 11450 2603 11452
rect 2357 11398 2359 11450
rect 2539 11398 2541 11450
rect 2295 11396 2301 11398
rect 2357 11396 2381 11398
rect 2437 11396 2461 11398
rect 2517 11396 2541 11398
rect 2597 11396 2603 11398
rect 2295 11387 2603 11396
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1872 10062 1900 10950
rect 2424 10810 2452 11018
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2502 10704 2558 10713
rect 2502 10639 2504 10648
rect 2556 10639 2558 10648
rect 2504 10610 2556 10616
rect 2792 10538 2820 10950
rect 2884 10792 2912 11494
rect 3252 11354 3280 11494
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3436 11098 3464 11494
rect 3608 11144 3660 11150
rect 3436 11092 3608 11098
rect 3436 11086 3660 11092
rect 3436 11070 3648 11086
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 2955 10908 3263 10917
rect 2955 10906 2961 10908
rect 3017 10906 3041 10908
rect 3097 10906 3121 10908
rect 3177 10906 3201 10908
rect 3257 10906 3263 10908
rect 3017 10854 3019 10906
rect 3199 10854 3201 10906
rect 2955 10852 2961 10854
rect 3017 10852 3041 10854
rect 3097 10852 3121 10854
rect 3177 10852 3201 10854
rect 3257 10852 3263 10854
rect 2955 10843 3263 10852
rect 2884 10764 3188 10792
rect 3056 10668 3108 10674
rect 2976 10628 3056 10656
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2295 10364 2603 10373
rect 2295 10362 2301 10364
rect 2357 10362 2381 10364
rect 2437 10362 2461 10364
rect 2517 10362 2541 10364
rect 2597 10362 2603 10364
rect 2357 10310 2359 10362
rect 2539 10310 2541 10362
rect 2295 10308 2301 10310
rect 2357 10308 2381 10310
rect 2437 10308 2461 10310
rect 2517 10308 2541 10310
rect 2597 10308 2603 10310
rect 2295 10299 2603 10308
rect 2792 10266 2820 10474
rect 2976 10266 3004 10628
rect 3056 10610 3108 10616
rect 3160 10606 3188 10764
rect 3344 10674 3372 10950
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 3068 10198 3096 10474
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 2504 10056 2556 10062
rect 2556 10004 2728 10010
rect 2504 9998 2728 10004
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 938 8871 994 8880
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1780 7818 1808 8434
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1872 7698 1900 9998
rect 2516 9994 2728 9998
rect 2516 9988 2740 9994
rect 2516 9982 2688 9988
rect 2688 9930 2740 9936
rect 2700 9654 2728 9930
rect 2955 9820 3263 9829
rect 2955 9818 2961 9820
rect 3017 9818 3041 9820
rect 3097 9818 3121 9820
rect 3177 9818 3201 9820
rect 3257 9818 3263 9820
rect 3017 9766 3019 9818
rect 3199 9766 3201 9818
rect 2955 9764 2961 9766
rect 3017 9764 3041 9766
rect 3097 9764 3121 9766
rect 3177 9764 3201 9766
rect 3257 9764 3263 9766
rect 2955 9755 3263 9764
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2295 9276 2603 9285
rect 2295 9274 2301 9276
rect 2357 9274 2381 9276
rect 2437 9274 2461 9276
rect 2517 9274 2541 9276
rect 2597 9274 2603 9276
rect 2357 9222 2359 9274
rect 2539 9222 2541 9274
rect 2295 9220 2301 9222
rect 2357 9220 2381 9222
rect 2437 9220 2461 9222
rect 2517 9220 2541 9222
rect 2597 9220 2603 9222
rect 2295 9211 2603 9220
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1780 7670 1900 7698
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 938 5536 994 5545
rect 938 5471 994 5480
rect 952 5302 980 5471
rect 1688 5302 1716 6734
rect 940 5296 992 5302
rect 940 5238 992 5244
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 952 2825 980 3402
rect 1596 3194 1624 4082
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 1780 2774 1808 7670
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1872 5914 1900 6802
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1964 5794 1992 7890
rect 2056 7886 2084 8842
rect 2700 8820 2728 9590
rect 3436 9586 3464 11070
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3528 10810 3556 10950
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3712 10674 3740 11834
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 4080 11354 4108 11766
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10674 3832 10950
rect 4540 10810 4568 11630
rect 4724 11014 4752 12242
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 5000 11898 5028 12106
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 5646 11996 5954 12005
rect 5646 11994 5652 11996
rect 5708 11994 5732 11996
rect 5788 11994 5812 11996
rect 5868 11994 5892 11996
rect 5948 11994 5954 11996
rect 5708 11942 5710 11994
rect 5890 11942 5892 11994
rect 5646 11940 5652 11942
rect 5708 11940 5732 11942
rect 5788 11940 5812 11942
rect 5868 11940 5892 11942
rect 5948 11940 5954 11942
rect 5646 11931 5954 11940
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4724 10674 4752 10950
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3792 10668 3844 10674
rect 4528 10668 4580 10674
rect 3792 10610 3844 10616
rect 4264 10628 4528 10656
rect 3528 10198 3556 10610
rect 3620 10266 3648 10610
rect 4160 10600 4212 10606
rect 4264 10588 4292 10628
rect 4528 10610 4580 10616
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4212 10560 4292 10588
rect 4160 10542 4212 10548
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3712 9994 3740 10202
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 2780 8832 2832 8838
rect 2700 8792 2780 8820
rect 2780 8774 2832 8780
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 2792 8514 2820 8774
rect 2884 8634 2912 8774
rect 2955 8732 3263 8741
rect 2955 8730 2961 8732
rect 3017 8730 3041 8732
rect 3097 8730 3121 8732
rect 3177 8730 3201 8732
rect 3257 8730 3263 8732
rect 3017 8678 3019 8730
rect 3199 8678 3201 8730
rect 2955 8676 2961 8678
rect 3017 8676 3041 8678
rect 3097 8676 3121 8678
rect 3177 8676 3201 8678
rect 3257 8676 3263 8678
rect 2955 8667 3263 8676
rect 3344 8634 3372 8774
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3436 8566 3464 9522
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9058 3648 9318
rect 3528 9030 3648 9058
rect 3528 8974 3556 9030
rect 3896 8974 3924 10066
rect 3988 9674 4016 10202
rect 4356 10146 4384 10474
rect 4540 10266 4568 10610
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4080 10118 4384 10146
rect 4080 10062 4108 10118
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 3988 9646 4200 9674
rect 4172 9178 4200 9646
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3424 8560 3476 8566
rect 2792 8486 3004 8514
rect 3424 8502 3476 8508
rect 2976 8430 3004 8486
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2240 8242 2268 8298
rect 2148 8214 2268 8242
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2056 6322 2084 6802
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1872 5766 1992 5794
rect 1872 3398 1900 5766
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1964 4826 1992 4966
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1964 4214 1992 4422
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 2056 3602 2084 5102
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2148 3534 2176 8214
rect 2295 8188 2603 8197
rect 2295 8186 2301 8188
rect 2357 8186 2381 8188
rect 2437 8186 2461 8188
rect 2517 8186 2541 8188
rect 2597 8186 2603 8188
rect 2357 8134 2359 8186
rect 2539 8134 2541 8186
rect 2295 8132 2301 8134
rect 2357 8132 2381 8134
rect 2437 8132 2461 8134
rect 2517 8132 2541 8134
rect 2597 8132 2603 8134
rect 2295 8123 2603 8132
rect 3528 7954 3556 8434
rect 3712 8362 3740 8910
rect 4264 8430 4292 9862
rect 4540 9674 4568 10202
rect 4816 10062 4844 10610
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4908 9926 4936 11630
rect 4986 11452 5294 11461
rect 4986 11450 4992 11452
rect 5048 11450 5072 11452
rect 5128 11450 5152 11452
rect 5208 11450 5232 11452
rect 5288 11450 5294 11452
rect 5048 11398 5050 11450
rect 5230 11398 5232 11450
rect 4986 11396 4992 11398
rect 5048 11396 5072 11398
rect 5128 11396 5152 11398
rect 5208 11396 5232 11398
rect 5288 11396 5294 11398
rect 4986 11387 5294 11396
rect 5368 10810 5396 11698
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11098 5488 11494
rect 5552 11218 5580 11630
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11354 5672 11494
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5460 11070 5580 11098
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5460 10713 5488 10950
rect 5446 10704 5502 10713
rect 5446 10639 5502 10648
rect 4986 10364 5294 10373
rect 4986 10362 4992 10364
rect 5048 10362 5072 10364
rect 5128 10362 5152 10364
rect 5208 10362 5232 10364
rect 5288 10362 5294 10364
rect 5048 10310 5050 10362
rect 5230 10310 5232 10362
rect 4986 10308 4992 10310
rect 5048 10308 5072 10310
rect 5128 10308 5152 10310
rect 5208 10308 5232 10310
rect 5288 10308 5294 10310
rect 4986 10299 5294 10308
rect 5460 10010 5488 10639
rect 5552 10130 5580 11070
rect 6012 11014 6040 11766
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6656 11150 6684 11494
rect 7677 11452 7985 11461
rect 7677 11450 7683 11452
rect 7739 11450 7763 11452
rect 7819 11450 7843 11452
rect 7899 11450 7923 11452
rect 7979 11450 7985 11452
rect 7739 11398 7741 11450
rect 7921 11398 7923 11450
rect 7677 11396 7683 11398
rect 7739 11396 7763 11398
rect 7819 11396 7843 11398
rect 7899 11396 7923 11398
rect 7979 11396 7985 11398
rect 7677 11387 7985 11396
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 5646 10908 5954 10917
rect 5646 10906 5652 10908
rect 5708 10906 5732 10908
rect 5788 10906 5812 10908
rect 5868 10906 5892 10908
rect 5948 10906 5954 10908
rect 5708 10854 5710 10906
rect 5890 10854 5892 10906
rect 5646 10852 5652 10854
rect 5708 10852 5732 10854
rect 5788 10852 5812 10854
rect 5868 10852 5892 10854
rect 5948 10852 5954 10854
rect 5646 10843 5954 10852
rect 6012 10810 6040 10950
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5908 10600 5960 10606
rect 6748 10554 6776 10950
rect 7024 10810 7052 11018
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 5908 10542 5960 10548
rect 5920 10266 5948 10542
rect 6656 10538 6776 10554
rect 6644 10532 6776 10538
rect 6696 10526 6776 10532
rect 6644 10474 6696 10480
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 6748 10130 6776 10406
rect 6840 10266 6868 10610
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 5460 9982 5580 10010
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4540 9646 4844 9674
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 2955 7644 3263 7653
rect 2955 7642 2961 7644
rect 3017 7642 3041 7644
rect 3097 7642 3121 7644
rect 3177 7642 3201 7644
rect 3257 7642 3263 7644
rect 3017 7590 3019 7642
rect 3199 7590 3201 7642
rect 2955 7588 2961 7590
rect 3017 7588 3041 7590
rect 3097 7588 3121 7590
rect 3177 7588 3201 7590
rect 3257 7588 3263 7590
rect 2955 7579 3263 7588
rect 3436 7546 3464 7822
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 2295 7100 2603 7109
rect 2295 7098 2301 7100
rect 2357 7098 2381 7100
rect 2437 7098 2461 7100
rect 2517 7098 2541 7100
rect 2597 7098 2603 7100
rect 2357 7046 2359 7098
rect 2539 7046 2541 7098
rect 2295 7044 2301 7046
rect 2357 7044 2381 7046
rect 2437 7044 2461 7046
rect 2517 7044 2541 7046
rect 2597 7044 2603 7046
rect 2295 7035 2603 7044
rect 3068 6798 3096 7482
rect 3528 7410 3556 7686
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3344 6662 3372 7278
rect 3436 6934 3464 7278
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3436 6798 3464 6870
rect 3528 6798 3556 7346
rect 3620 7002 3648 7822
rect 3804 7478 3832 8230
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 2240 6458 2268 6598
rect 2955 6556 3263 6565
rect 2955 6554 2961 6556
rect 3017 6554 3041 6556
rect 3097 6554 3121 6556
rect 3177 6554 3201 6556
rect 3257 6554 3263 6556
rect 3017 6502 3019 6554
rect 3199 6502 3201 6554
rect 2955 6500 2961 6502
rect 3017 6500 3041 6502
rect 3097 6500 3121 6502
rect 3177 6500 3201 6502
rect 3257 6500 3263 6502
rect 2955 6491 3263 6500
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2295 6012 2603 6021
rect 2295 6010 2301 6012
rect 2357 6010 2381 6012
rect 2437 6010 2461 6012
rect 2517 6010 2541 6012
rect 2597 6010 2603 6012
rect 2357 5958 2359 6010
rect 2539 5958 2541 6010
rect 2295 5956 2301 5958
rect 2357 5956 2381 5958
rect 2437 5956 2461 5958
rect 2517 5956 2541 5958
rect 2597 5956 2603 5958
rect 2295 5947 2603 5956
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2608 5250 2636 5646
rect 2700 5370 2728 6122
rect 2976 5574 3004 6122
rect 3344 5778 3372 6598
rect 3528 6458 3556 6734
rect 3896 6730 3924 7278
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3884 6724 3936 6730
rect 3884 6666 3936 6672
rect 3896 6458 3924 6666
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3896 5914 3924 6190
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 4172 5778 4200 7142
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 2955 5468 3263 5477
rect 2955 5466 2961 5468
rect 3017 5466 3041 5468
rect 3097 5466 3121 5468
rect 3177 5466 3201 5468
rect 3257 5466 3263 5468
rect 3017 5414 3019 5466
rect 3199 5414 3201 5466
rect 2955 5412 2961 5414
rect 3017 5412 3041 5414
rect 3097 5412 3121 5414
rect 3177 5412 3201 5414
rect 3257 5412 3263 5414
rect 2955 5403 3263 5412
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 3332 5296 3384 5302
rect 2608 5222 2728 5250
rect 3332 5238 3384 5244
rect 2295 4924 2603 4933
rect 2295 4922 2301 4924
rect 2357 4922 2381 4924
rect 2437 4922 2461 4924
rect 2517 4922 2541 4924
rect 2597 4922 2603 4924
rect 2357 4870 2359 4922
rect 2539 4870 2541 4922
rect 2295 4868 2301 4870
rect 2357 4868 2381 4870
rect 2437 4868 2461 4870
rect 2517 4868 2541 4870
rect 2597 4868 2603 4870
rect 2295 4859 2603 4868
rect 2700 4282 2728 5222
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2295 3836 2603 3845
rect 2295 3834 2301 3836
rect 2357 3834 2381 3836
rect 2437 3834 2461 3836
rect 2517 3834 2541 3836
rect 2597 3834 2603 3836
rect 2357 3782 2359 3834
rect 2539 3782 2541 3834
rect 2295 3780 2301 3782
rect 2357 3780 2381 3782
rect 2437 3780 2461 3782
rect 2517 3780 2541 3782
rect 2597 3780 2603 3782
rect 2295 3771 2603 3780
rect 2700 3670 2728 4218
rect 2884 4010 2912 4966
rect 2955 4380 3263 4389
rect 2955 4378 2961 4380
rect 3017 4378 3041 4380
rect 3097 4378 3121 4380
rect 3177 4378 3201 4380
rect 3257 4378 3263 4380
rect 3017 4326 3019 4378
rect 3199 4326 3201 4378
rect 2955 4324 2961 4326
rect 3017 4324 3041 4326
rect 3097 4324 3121 4326
rect 3177 4324 3201 4326
rect 3257 4324 3263 4326
rect 2955 4315 3263 4324
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 3344 3942 3372 5238
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3528 3738 3556 4150
rect 3712 4146 3740 5510
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3804 4078 3832 4422
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 4080 3534 4108 4150
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2332 2854 2360 3334
rect 2792 3108 2820 3334
rect 2955 3292 3263 3301
rect 2955 3290 2961 3292
rect 3017 3290 3041 3292
rect 3097 3290 3121 3292
rect 3177 3290 3201 3292
rect 3257 3290 3263 3292
rect 3017 3238 3019 3290
rect 3199 3238 3201 3290
rect 2955 3236 2961 3238
rect 3017 3236 3041 3238
rect 3097 3236 3121 3238
rect 3177 3236 3201 3238
rect 3257 3236 3263 3238
rect 2955 3227 3263 3236
rect 4080 3126 4108 3470
rect 2700 3080 2820 3108
rect 4068 3120 4120 3126
rect 2700 2990 2728 3080
rect 4068 3062 4120 3068
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 1780 2746 1900 2774
rect 1872 2446 1900 2746
rect 2295 2748 2603 2757
rect 2295 2746 2301 2748
rect 2357 2746 2381 2748
rect 2437 2746 2461 2748
rect 2517 2746 2541 2748
rect 2597 2746 2603 2748
rect 2357 2694 2359 2746
rect 2539 2694 2541 2746
rect 2295 2692 2301 2694
rect 2357 2692 2381 2694
rect 2437 2692 2461 2694
rect 2517 2692 2541 2694
rect 2597 2692 2603 2694
rect 2295 2683 2603 2692
rect 4172 2514 4200 4218
rect 4264 4078 4292 8366
rect 4540 6458 4568 8842
rect 4632 8634 4660 8842
rect 4724 8634 4752 9114
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4632 7342 4660 8366
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4356 5914 4384 6258
rect 4448 6118 4476 6326
rect 4816 6202 4844 9646
rect 4724 6174 4844 6202
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4448 5166 4476 6054
rect 4724 5914 4752 6174
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4816 5710 4844 6054
rect 4908 5778 4936 9862
rect 5552 9654 5580 9982
rect 6932 9926 6960 10746
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7116 10198 7144 10542
rect 7392 10266 7420 10610
rect 7677 10364 7985 10373
rect 7677 10362 7683 10364
rect 7739 10362 7763 10364
rect 7819 10362 7843 10364
rect 7899 10362 7923 10364
rect 7979 10362 7985 10364
rect 7739 10310 7741 10362
rect 7921 10310 7923 10362
rect 7677 10308 7683 10310
rect 7739 10308 7763 10310
rect 7819 10308 7843 10310
rect 7899 10308 7923 10310
rect 7979 10308 7985 10310
rect 7677 10299 7985 10308
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 5646 9820 5954 9829
rect 5646 9818 5652 9820
rect 5708 9818 5732 9820
rect 5788 9818 5812 9820
rect 5868 9818 5892 9820
rect 5948 9818 5954 9820
rect 5708 9766 5710 9818
rect 5890 9766 5892 9818
rect 5646 9764 5652 9766
rect 5708 9764 5732 9766
rect 5788 9764 5812 9766
rect 5868 9764 5892 9766
rect 5948 9764 5954 9766
rect 5646 9755 5954 9764
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 4986 9276 5294 9285
rect 4986 9274 4992 9276
rect 5048 9274 5072 9276
rect 5128 9274 5152 9276
rect 5208 9274 5232 9276
rect 5288 9274 5294 9276
rect 5048 9222 5050 9274
rect 5230 9222 5232 9274
rect 4986 9220 4992 9222
rect 5048 9220 5072 9222
rect 5128 9220 5152 9222
rect 5208 9220 5232 9222
rect 5288 9220 5294 9222
rect 4986 9211 5294 9220
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 8634 5212 8842
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 4986 8188 5294 8197
rect 4986 8186 4992 8188
rect 5048 8186 5072 8188
rect 5128 8186 5152 8188
rect 5208 8186 5232 8188
rect 5288 8186 5294 8188
rect 5048 8134 5050 8186
rect 5230 8134 5232 8186
rect 4986 8132 4992 8134
rect 5048 8132 5072 8134
rect 5128 8132 5152 8134
rect 5208 8132 5232 8134
rect 5288 8132 5294 8134
rect 4986 8123 5294 8132
rect 4986 7100 5294 7109
rect 4986 7098 4992 7100
rect 5048 7098 5072 7100
rect 5128 7098 5152 7100
rect 5208 7098 5232 7100
rect 5288 7098 5294 7100
rect 5048 7046 5050 7098
rect 5230 7046 5232 7098
rect 4986 7044 4992 7046
rect 5048 7044 5072 7046
rect 5128 7044 5152 7046
rect 5208 7044 5232 7046
rect 5288 7044 5294 7046
rect 4986 7035 5294 7044
rect 5368 6798 5396 9114
rect 7024 9042 7052 9590
rect 7677 9276 7985 9285
rect 7677 9274 7683 9276
rect 7739 9274 7763 9276
rect 7819 9274 7843 9276
rect 7899 9274 7923 9276
rect 7979 9274 7985 9276
rect 7739 9222 7741 9274
rect 7921 9222 7923 9274
rect 7677 9220 7683 9222
rect 7739 9220 7763 9222
rect 7819 9220 7843 9222
rect 7899 9220 7923 9222
rect 7979 9220 7985 9222
rect 7677 9211 7985 9220
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 5646 8732 5954 8741
rect 5646 8730 5652 8732
rect 5708 8730 5732 8732
rect 5788 8730 5812 8732
rect 5868 8730 5892 8732
rect 5948 8730 5954 8732
rect 5708 8678 5710 8730
rect 5890 8678 5892 8730
rect 5646 8676 5652 8678
rect 5708 8676 5732 8678
rect 5788 8676 5812 8678
rect 5868 8676 5892 8678
rect 5948 8676 5954 8678
rect 5646 8667 5954 8676
rect 6196 8634 6224 8842
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6380 8498 6408 8978
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 5646 7644 5954 7653
rect 5646 7642 5652 7644
rect 5708 7642 5732 7644
rect 5788 7642 5812 7644
rect 5868 7642 5892 7644
rect 5948 7642 5954 7644
rect 5708 7590 5710 7642
rect 5890 7590 5892 7642
rect 5646 7588 5652 7590
rect 5708 7588 5732 7590
rect 5788 7588 5812 7590
rect 5868 7588 5892 7590
rect 5948 7588 5954 7590
rect 5646 7579 5954 7588
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5184 6458 5212 6666
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5092 6186 5120 6394
rect 5368 6322 5396 6734
rect 5552 6322 5580 7142
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5646 6556 5954 6565
rect 5646 6554 5652 6556
rect 5708 6554 5732 6556
rect 5788 6554 5812 6556
rect 5868 6554 5892 6556
rect 5948 6554 5954 6556
rect 5708 6502 5710 6554
rect 5890 6502 5892 6554
rect 5646 6500 5652 6502
rect 5708 6500 5732 6502
rect 5788 6500 5812 6502
rect 5868 6500 5892 6502
rect 5948 6500 5954 6502
rect 5646 6491 5954 6500
rect 6012 6458 6040 6598
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5276 6100 5304 6258
rect 5540 6112 5592 6118
rect 5276 6072 5396 6100
rect 4986 6012 5294 6021
rect 4986 6010 4992 6012
rect 5048 6010 5072 6012
rect 5128 6010 5152 6012
rect 5208 6010 5232 6012
rect 5288 6010 5294 6012
rect 5048 5958 5050 6010
rect 5230 5958 5232 6010
rect 4986 5956 4992 5958
rect 5048 5956 5072 5958
rect 5128 5956 5152 5958
rect 5208 5956 5232 5958
rect 5288 5956 5294 5958
rect 4986 5947 5294 5956
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4448 4690 4476 5102
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4540 3126 4568 5510
rect 4724 5370 4752 5646
rect 4908 5370 4936 5714
rect 5092 5710 5120 5850
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4908 4622 4936 5306
rect 5368 5234 5396 6072
rect 5540 6054 5592 6060
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5552 5710 5580 6054
rect 5644 5778 5672 6054
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5540 5704 5592 5710
rect 5460 5652 5540 5658
rect 5460 5646 5592 5652
rect 5460 5630 5580 5646
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 4986 4924 5294 4933
rect 4986 4922 4992 4924
rect 5048 4922 5072 4924
rect 5128 4922 5152 4924
rect 5208 4922 5232 4924
rect 5288 4922 5294 4924
rect 5048 4870 5050 4922
rect 5230 4870 5232 4922
rect 4986 4868 4992 4870
rect 5048 4868 5072 4870
rect 5128 4868 5152 4870
rect 5208 4868 5232 4870
rect 5288 4868 5294 4870
rect 4986 4859 5294 4868
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 5460 4282 5488 5630
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 4826 5580 5510
rect 5646 5468 5954 5477
rect 5646 5466 5652 5468
rect 5708 5466 5732 5468
rect 5788 5466 5812 5468
rect 5868 5466 5892 5468
rect 5948 5466 5954 5468
rect 5708 5414 5710 5466
rect 5890 5414 5892 5466
rect 5646 5412 5652 5414
rect 5708 5412 5732 5414
rect 5788 5412 5812 5414
rect 5868 5412 5892 5414
rect 5948 5412 5954 5414
rect 5646 5403 5954 5412
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5646 4380 5954 4389
rect 5646 4378 5652 4380
rect 5708 4378 5732 4380
rect 5788 4378 5812 4380
rect 5868 4378 5892 4380
rect 5948 4378 5954 4380
rect 5708 4326 5710 4378
rect 5890 4326 5892 4378
rect 5646 4324 5652 4326
rect 5708 4324 5732 4326
rect 5788 4324 5812 4326
rect 5868 4324 5892 4326
rect 5948 4324 5954 4326
rect 5646 4315 5954 4324
rect 6104 4282 6132 8366
rect 6380 8090 6408 8434
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6274 6760 6330 6769
rect 6274 6695 6330 6704
rect 6288 6662 6316 6695
rect 6564 6662 6592 8502
rect 7024 8430 7052 8978
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8566 7144 8774
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 8036 8362 8064 12038
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7677 8188 7985 8197
rect 7677 8186 7683 8188
rect 7739 8186 7763 8188
rect 7819 8186 7843 8188
rect 7899 8186 7923 8188
rect 7979 8186 7985 8188
rect 7739 8134 7741 8186
rect 7921 8134 7923 8186
rect 7677 8132 7683 8134
rect 7739 8132 7763 8134
rect 7819 8132 7843 8134
rect 7899 8132 7923 8134
rect 7979 8132 7985 8134
rect 7677 8123 7985 8132
rect 8036 7954 8064 8298
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 7206 6960 7754
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 7041 6960 7142
rect 6918 7032 6974 7041
rect 6828 6996 6880 7002
rect 6918 6967 6974 6976
rect 6828 6938 6880 6944
rect 6840 6798 6868 6938
rect 7300 6798 7328 7686
rect 7677 7100 7985 7109
rect 7677 7098 7683 7100
rect 7739 7098 7763 7100
rect 7819 7098 7843 7100
rect 7899 7098 7923 7100
rect 7979 7098 7985 7100
rect 7739 7046 7741 7098
rect 7921 7046 7923 7098
rect 7677 7044 7683 7046
rect 7739 7044 7763 7046
rect 7819 7044 7843 7046
rect 7899 7044 7923 7046
rect 7979 7044 7985 7046
rect 7677 7035 7985 7044
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7562 6760 7618 6769
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6288 6390 6316 6598
rect 6276 6384 6328 6390
rect 6932 6361 6960 6734
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6474 7328 6598
rect 7024 6458 7328 6474
rect 7012 6452 7328 6458
rect 7064 6446 7328 6452
rect 7012 6394 7064 6400
rect 6276 6326 6328 6332
rect 6918 6352 6974 6361
rect 7392 6338 7420 6734
rect 7472 6724 7524 6730
rect 7562 6695 7618 6704
rect 7472 6666 7524 6672
rect 7484 6440 7512 6666
rect 7576 6662 7604 6695
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7564 6452 7616 6458
rect 7484 6412 7564 6440
rect 7564 6394 7616 6400
rect 6918 6287 6974 6296
rect 7300 6310 7420 6338
rect 8036 6322 8064 7890
rect 8128 6338 8156 12106
rect 8337 11996 8645 12005
rect 8337 11994 8343 11996
rect 8399 11994 8423 11996
rect 8479 11994 8503 11996
rect 8559 11994 8583 11996
rect 8639 11994 8645 11996
rect 8399 11942 8401 11994
rect 8581 11942 8583 11994
rect 8337 11940 8343 11942
rect 8399 11940 8423 11942
rect 8479 11940 8503 11942
rect 8559 11940 8583 11942
rect 8639 11940 8645 11942
rect 8337 11931 8645 11940
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8312 11150 8340 11698
rect 8680 11354 8708 12174
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9048 11898 9076 12038
rect 10152 11898 10180 12242
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11028 11996 11336 12005
rect 11028 11994 11034 11996
rect 11090 11994 11114 11996
rect 11170 11994 11194 11996
rect 11250 11994 11274 11996
rect 11330 11994 11336 11996
rect 11090 11942 11092 11994
rect 11272 11942 11274 11994
rect 11028 11940 11034 11942
rect 11090 11940 11114 11942
rect 11170 11940 11194 11942
rect 11250 11940 11274 11942
rect 11330 11940 11336 11942
rect 11028 11931 11336 11940
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8337 10908 8645 10917
rect 8337 10906 8343 10908
rect 8399 10906 8423 10908
rect 8479 10906 8503 10908
rect 8559 10906 8583 10908
rect 8639 10906 8645 10908
rect 8399 10854 8401 10906
rect 8581 10854 8583 10906
rect 8337 10852 8343 10854
rect 8399 10852 8423 10854
rect 8479 10852 8503 10854
rect 8559 10852 8583 10854
rect 8639 10852 8645 10854
rect 8337 10843 8645 10852
rect 8680 10674 8708 11290
rect 8772 11014 8800 11494
rect 8864 11218 8892 11494
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8220 10130 8248 10474
rect 8312 10470 8340 10610
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8312 10062 8340 10406
rect 8404 10198 8432 10610
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8680 9926 8708 10610
rect 8772 10130 8800 10950
rect 8956 10742 8984 10950
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 9600 10606 9628 11494
rect 9784 11354 9812 11766
rect 10368 11452 10676 11461
rect 10368 11450 10374 11452
rect 10430 11450 10454 11452
rect 10510 11450 10534 11452
rect 10590 11450 10614 11452
rect 10670 11450 10676 11452
rect 10430 11398 10432 11450
rect 10612 11398 10614 11450
rect 10368 11396 10374 11398
rect 10430 11396 10454 11398
rect 10510 11396 10534 11398
rect 10590 11396 10614 11398
rect 10670 11396 10676 11398
rect 10368 11387 10676 11396
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8337 9820 8645 9829
rect 8337 9818 8343 9820
rect 8399 9818 8423 9820
rect 8479 9818 8503 9820
rect 8559 9818 8583 9820
rect 8639 9818 8645 9820
rect 8399 9766 8401 9818
rect 8581 9766 8583 9818
rect 8337 9764 8343 9766
rect 8399 9764 8423 9766
rect 8479 9764 8503 9766
rect 8559 9764 8583 9766
rect 8639 9764 8645 9766
rect 8337 9755 8645 9764
rect 9324 9654 9352 10134
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8772 9042 8800 9318
rect 8864 9178 8892 9386
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8956 9110 8984 9454
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8337 8732 8645 8741
rect 8337 8730 8343 8732
rect 8399 8730 8423 8732
rect 8479 8730 8503 8732
rect 8559 8730 8583 8732
rect 8639 8730 8645 8732
rect 8399 8678 8401 8730
rect 8581 8678 8583 8730
rect 8337 8676 8343 8678
rect 8399 8676 8423 8678
rect 8479 8676 8503 8678
rect 8559 8676 8583 8678
rect 8639 8676 8645 8678
rect 8337 8667 8645 8676
rect 8864 8566 8892 8910
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8956 8566 8984 8774
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9048 8090 9076 8434
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8337 7644 8645 7653
rect 8337 7642 8343 7644
rect 8399 7642 8423 7644
rect 8479 7642 8503 7644
rect 8559 7642 8583 7644
rect 8639 7642 8645 7644
rect 8399 7590 8401 7642
rect 8581 7590 8583 7642
rect 8337 7588 8343 7590
rect 8399 7588 8423 7590
rect 8479 7588 8503 7590
rect 8559 7588 8583 7590
rect 8639 7588 8645 7590
rect 8337 7579 8645 7588
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8220 7041 8248 7346
rect 8206 7032 8262 7041
rect 8206 6967 8262 6976
rect 8337 6556 8645 6565
rect 8337 6554 8343 6556
rect 8399 6554 8423 6556
rect 8479 6554 8503 6556
rect 8559 6554 8583 6556
rect 8639 6554 8645 6556
rect 8399 6502 8401 6554
rect 8581 6502 8583 6554
rect 8337 6500 8343 6502
rect 8399 6500 8423 6502
rect 8479 6500 8503 6502
rect 8559 6500 8583 6502
rect 8639 6500 8645 6502
rect 8337 6491 8645 6500
rect 8484 6384 8536 6390
rect 8128 6322 8340 6338
rect 8484 6326 8536 6332
rect 8024 6316 8076 6322
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6840 5846 6868 6190
rect 6932 5914 6960 6287
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6288 4622 6316 5646
rect 6840 5234 6868 5782
rect 7024 5352 7052 6054
rect 7116 5642 7144 6190
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 7024 5324 7144 5352
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6840 4690 6868 5170
rect 7116 4758 7144 5324
rect 7300 5234 7328 6310
rect 8024 6258 8076 6264
rect 8128 6316 8352 6322
rect 8128 6310 8300 6316
rect 7677 6012 7985 6021
rect 7677 6010 7683 6012
rect 7739 6010 7763 6012
rect 7819 6010 7843 6012
rect 7899 6010 7923 6012
rect 7979 6010 7985 6012
rect 7739 5958 7741 6010
rect 7921 5958 7923 6010
rect 7677 5956 7683 5958
rect 7739 5956 7763 5958
rect 7819 5956 7843 5958
rect 7899 5956 7923 5958
rect 7979 5956 7985 5958
rect 7677 5947 7985 5956
rect 8036 5692 8064 6258
rect 8128 5914 8156 6310
rect 8300 6258 8352 6264
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8220 5710 8248 6190
rect 8496 6118 8524 6326
rect 8680 6254 8708 7890
rect 9140 7886 9168 9590
rect 9508 9110 9536 10406
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9416 8974 9444 9046
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8680 5914 8708 6190
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8116 5704 8168 5710
rect 8036 5664 8116 5692
rect 8116 5646 8168 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8588 5658 8616 5714
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6182 4040 6238 4049
rect 5540 4004 5592 4010
rect 6182 3975 6238 3984
rect 5540 3946 5592 3952
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 4986 3836 5294 3845
rect 4986 3834 4992 3836
rect 5048 3834 5072 3836
rect 5128 3834 5152 3836
rect 5208 3834 5232 3836
rect 5288 3834 5294 3836
rect 5048 3782 5050 3834
rect 5230 3782 5232 3834
rect 4986 3780 4992 3782
rect 5048 3780 5072 3782
rect 5128 3780 5152 3782
rect 5208 3780 5232 3782
rect 5288 3780 5294 3782
rect 4986 3771 5294 3780
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4816 3194 4844 3538
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5460 3126 5488 3878
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5552 2774 5580 3946
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5646 3292 5954 3301
rect 5646 3290 5652 3292
rect 5708 3290 5732 3292
rect 5788 3290 5812 3292
rect 5868 3290 5892 3292
rect 5948 3290 5954 3292
rect 5708 3238 5710 3290
rect 5890 3238 5892 3290
rect 5646 3236 5652 3238
rect 5708 3236 5732 3238
rect 5788 3236 5812 3238
rect 5868 3236 5892 3238
rect 5948 3236 5954 3238
rect 5646 3227 5954 3236
rect 4986 2748 5294 2757
rect 4986 2746 4992 2748
rect 5048 2746 5072 2748
rect 5128 2746 5152 2748
rect 5208 2746 5232 2748
rect 5288 2746 5294 2748
rect 5552 2746 5764 2774
rect 5048 2694 5050 2746
rect 5230 2694 5232 2746
rect 4986 2692 4992 2694
rect 5048 2692 5072 2694
rect 5128 2692 5152 2694
rect 5208 2692 5232 2694
rect 5288 2692 5294 2694
rect 4986 2683 5294 2692
rect 5736 2514 5764 2746
rect 6012 2514 6040 3538
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 5460 2378 5672 2394
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 5460 2372 5684 2378
rect 5460 2366 5632 2372
rect 32 800 60 2314
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 800 2636 2246
rect 2955 2204 3263 2213
rect 2955 2202 2961 2204
rect 3017 2202 3041 2204
rect 3097 2202 3121 2204
rect 3177 2202 3201 2204
rect 3257 2202 3263 2204
rect 3017 2150 3019 2202
rect 3199 2150 3201 2202
rect 2955 2148 2961 2150
rect 3017 2148 3041 2150
rect 3097 2148 3121 2150
rect 3177 2148 3201 2150
rect 3257 2148 3263 2150
rect 2955 2139 3263 2148
rect 5184 870 5304 898
rect 5184 800 5212 870
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 5276 762 5304 870
rect 5460 762 5488 2366
rect 5632 2314 5684 2320
rect 6104 2310 6132 3878
rect 6196 3534 6224 3975
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6184 2984 6236 2990
rect 6288 2972 6316 4558
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6236 2944 6316 2972
rect 6184 2926 6236 2932
rect 6196 2582 6224 2926
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 6472 2446 6500 4082
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6564 3194 6592 3402
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 7208 3126 7236 4422
rect 7300 3738 7328 5170
rect 7677 4924 7985 4933
rect 7677 4922 7683 4924
rect 7739 4922 7763 4924
rect 7819 4922 7843 4924
rect 7899 4922 7923 4924
rect 7979 4922 7985 4924
rect 7739 4870 7741 4922
rect 7921 4870 7923 4922
rect 7677 4868 7683 4870
rect 7739 4868 7763 4870
rect 7819 4868 7843 4870
rect 7899 4868 7923 4870
rect 7979 4868 7985 4870
rect 7677 4859 7985 4868
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7300 2650 7328 3402
rect 7576 3194 7604 4422
rect 7677 3836 7985 3845
rect 7677 3834 7683 3836
rect 7739 3834 7763 3836
rect 7819 3834 7843 3836
rect 7899 3834 7923 3836
rect 7979 3834 7985 3836
rect 7739 3782 7741 3834
rect 7921 3782 7923 3834
rect 7677 3780 7683 3782
rect 7739 3780 7763 3782
rect 7819 3780 7843 3782
rect 7899 3780 7923 3782
rect 7979 3780 7985 3782
rect 7677 3771 7985 3780
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7668 2990 7696 3674
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7760 3058 7788 3538
rect 8220 3466 8248 5646
rect 8588 5630 8708 5658
rect 8337 5468 8645 5477
rect 8337 5466 8343 5468
rect 8399 5466 8423 5468
rect 8479 5466 8503 5468
rect 8559 5466 8583 5468
rect 8639 5466 8645 5468
rect 8399 5414 8401 5466
rect 8581 5414 8583 5466
rect 8337 5412 8343 5414
rect 8399 5412 8423 5414
rect 8479 5412 8503 5414
rect 8559 5412 8583 5414
rect 8639 5412 8645 5414
rect 8337 5403 8645 5412
rect 8680 4622 8708 5630
rect 8772 5234 8800 6734
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8864 5778 8892 6598
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8956 5914 8984 6394
rect 9034 6352 9090 6361
rect 9034 6287 9090 6296
rect 9048 6254 9076 6287
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8772 4758 8800 5170
rect 8760 4752 8812 4758
rect 8760 4694 8812 4700
rect 8864 4690 8892 5578
rect 8956 5574 8984 5850
rect 9048 5778 9076 6054
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 9048 5302 9076 5714
rect 9140 5370 9168 6734
rect 9232 5914 9260 6734
rect 9416 6662 9444 8910
rect 9600 8498 9628 10542
rect 9692 10010 9720 11086
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9784 10130 9812 11018
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10742 9996 10950
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 10152 10266 10180 11086
rect 11028 10908 11336 10917
rect 11028 10906 11034 10908
rect 11090 10906 11114 10908
rect 11170 10906 11194 10908
rect 11250 10906 11274 10908
rect 11330 10906 11336 10908
rect 11090 10854 11092 10906
rect 11272 10854 11274 10906
rect 11028 10852 11034 10854
rect 11090 10852 11114 10854
rect 11170 10852 11194 10854
rect 11250 10852 11274 10854
rect 11330 10852 11336 10854
rect 11028 10843 11336 10852
rect 11440 10810 11468 12174
rect 12912 11898 12940 14346
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10368 10364 10676 10373
rect 10368 10362 10374 10364
rect 10430 10362 10454 10364
rect 10510 10362 10534 10364
rect 10590 10362 10614 10364
rect 10670 10362 10676 10364
rect 10430 10310 10432 10362
rect 10612 10310 10614 10362
rect 10368 10308 10374 10310
rect 10430 10308 10454 10310
rect 10510 10308 10534 10310
rect 10590 10308 10614 10310
rect 10670 10308 10676 10310
rect 10368 10299 10676 10308
rect 10888 10266 10916 10678
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9692 9982 9812 10010
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9518 9720 9862
rect 9784 9722 9812 9982
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 9178 9720 9318
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 9042 9812 9522
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9692 7954 9720 8026
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 6934 9720 7890
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9508 6458 9536 6666
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9324 6118 9352 6258
rect 9496 6248 9548 6254
rect 9416 6208 9496 6236
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9324 5778 9352 6054
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9416 5658 9444 6208
rect 9496 6190 9548 6196
rect 9600 5778 9628 6802
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9784 6254 9812 8978
rect 9876 8650 9904 10134
rect 11440 10062 11468 10746
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9968 9722 9996 9930
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9968 9602 9996 9658
rect 9968 9574 10088 9602
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 8838 9996 9318
rect 10060 9178 10088 9574
rect 10368 9276 10676 9285
rect 10368 9274 10374 9276
rect 10430 9274 10454 9276
rect 10510 9274 10534 9276
rect 10590 9274 10614 9276
rect 10670 9274 10676 9276
rect 10430 9222 10432 9274
rect 10612 9222 10614 9274
rect 10368 9220 10374 9222
rect 10430 9220 10454 9222
rect 10510 9220 10534 9222
rect 10590 9220 10614 9222
rect 10670 9220 10676 9222
rect 10368 9211 10676 9220
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9876 8622 9996 8650
rect 10152 8634 10180 8842
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9876 7954 9904 8230
rect 9968 8090 9996 8622
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10244 8090 10272 8366
rect 10368 8188 10676 8197
rect 10368 8186 10374 8188
rect 10430 8186 10454 8188
rect 10510 8186 10534 8188
rect 10590 8186 10614 8188
rect 10670 8186 10676 8188
rect 10430 8134 10432 8186
rect 10612 8134 10614 8186
rect 10368 8132 10374 8134
rect 10430 8132 10454 8134
rect 10510 8132 10534 8134
rect 10590 8132 10614 8134
rect 10670 8132 10676 8134
rect 10368 8123 10676 8132
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10704 8022 10732 9998
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11028 9820 11336 9829
rect 11028 9818 11034 9820
rect 11090 9818 11114 9820
rect 11170 9818 11194 9820
rect 11250 9818 11274 9820
rect 11330 9818 11336 9820
rect 11090 9766 11092 9818
rect 11272 9766 11274 9818
rect 11028 9764 11034 9766
rect 11090 9764 11114 9766
rect 11170 9764 11194 9766
rect 11250 9764 11274 9766
rect 11330 9764 11336 9766
rect 11028 9755 11336 9764
rect 11532 9382 11560 9930
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12084 9625 12112 9658
rect 12070 9616 12126 9625
rect 12070 9551 12126 9560
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11028 8732 11336 8741
rect 11028 8730 11034 8732
rect 11090 8730 11114 8732
rect 11170 8730 11194 8732
rect 11250 8730 11274 8732
rect 11330 8730 11336 8732
rect 11090 8678 11092 8730
rect 11272 8678 11274 8730
rect 11028 8676 11034 8678
rect 11090 8676 11114 8678
rect 11170 8676 11194 8678
rect 11250 8676 11274 8678
rect 11330 8676 11336 8678
rect 11028 8667 11336 8676
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 10368 7100 10676 7109
rect 10368 7098 10374 7100
rect 10430 7098 10454 7100
rect 10510 7098 10534 7100
rect 10590 7098 10614 7100
rect 10670 7098 10676 7100
rect 10430 7046 10432 7098
rect 10612 7046 10614 7098
rect 10368 7044 10374 7046
rect 10430 7044 10454 7046
rect 10510 7044 10534 7046
rect 10590 7044 10614 7046
rect 10670 7044 10676 7046
rect 10368 7035 10676 7044
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9324 5630 9444 5658
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9232 4826 9260 4966
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 8337 4380 8645 4389
rect 8337 4378 8343 4380
rect 8399 4378 8423 4380
rect 8479 4378 8503 4380
rect 8559 4378 8583 4380
rect 8639 4378 8645 4380
rect 8399 4326 8401 4378
rect 8581 4326 8583 4378
rect 8337 4324 8343 4326
rect 8399 4324 8423 4326
rect 8479 4324 8503 4326
rect 8559 4324 8583 4326
rect 8639 4324 8645 4326
rect 8337 4315 8645 4324
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7852 3194 7880 3334
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 8128 2990 8156 3334
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 7677 2748 7985 2757
rect 7677 2746 7683 2748
rect 7739 2746 7763 2748
rect 7819 2746 7843 2748
rect 7899 2746 7923 2748
rect 7979 2746 7985 2748
rect 7739 2694 7741 2746
rect 7921 2694 7923 2746
rect 7677 2692 7683 2694
rect 7739 2692 7763 2694
rect 7819 2692 7843 2694
rect 7899 2692 7923 2694
rect 7979 2692 7985 2694
rect 7677 2683 7985 2692
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 8220 2446 8248 3402
rect 8337 3292 8645 3301
rect 8337 3290 8343 3292
rect 8399 3290 8423 3292
rect 8479 3290 8503 3292
rect 8559 3290 8583 3292
rect 8639 3290 8645 3292
rect 8399 3238 8401 3290
rect 8581 3238 8583 3290
rect 8337 3236 8343 3238
rect 8399 3236 8423 3238
rect 8479 3236 8503 3238
rect 8559 3236 8583 3238
rect 8639 3236 8645 3238
rect 8337 3227 8645 3236
rect 8772 3126 8800 3878
rect 9140 3534 9168 4558
rect 9324 3670 9352 5630
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5370 9444 5510
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9508 5234 9536 5646
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9600 5098 9628 5714
rect 9784 5642 9812 6190
rect 9876 5914 9904 6734
rect 10368 6012 10676 6021
rect 10368 6010 10374 6012
rect 10430 6010 10454 6012
rect 10510 6010 10534 6012
rect 10590 6010 10614 6012
rect 10670 6010 10676 6012
rect 10430 5958 10432 6010
rect 10612 5958 10614 6010
rect 10368 5956 10374 5958
rect 10430 5956 10454 5958
rect 10510 5956 10534 5958
rect 10590 5956 10614 5958
rect 10670 5956 10676 5958
rect 10368 5947 10676 5956
rect 10704 5914 10732 7958
rect 10796 7750 10824 8570
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10888 8090 10916 8502
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9588 5092 9640 5098
rect 9588 5034 9640 5040
rect 10060 4690 10088 5510
rect 10368 4924 10676 4933
rect 10368 4922 10374 4924
rect 10430 4922 10454 4924
rect 10510 4922 10534 4924
rect 10590 4922 10614 4924
rect 10670 4922 10676 4924
rect 10430 4870 10432 4922
rect 10612 4870 10614 4922
rect 10368 4868 10374 4870
rect 10430 4868 10454 4870
rect 10510 4868 10534 4870
rect 10590 4868 10614 4870
rect 10670 4868 10676 4870
rect 10368 4859 10676 4868
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 9600 3602 9628 4422
rect 10704 4146 10732 5850
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10368 3836 10676 3845
rect 10368 3834 10374 3836
rect 10430 3834 10454 3836
rect 10510 3834 10534 3836
rect 10590 3834 10614 3836
rect 10670 3834 10676 3836
rect 10430 3782 10432 3834
rect 10612 3782 10614 3834
rect 10368 3780 10374 3782
rect 10430 3780 10454 3782
rect 10510 3780 10534 3782
rect 10590 3780 10614 3782
rect 10670 3780 10676 3782
rect 10368 3771 10676 3780
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9324 3194 9352 3470
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 9324 2774 9352 3130
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 9324 2746 9536 2774
rect 9508 2446 9536 2746
rect 10368 2748 10676 2757
rect 10368 2746 10374 2748
rect 10430 2746 10454 2748
rect 10510 2746 10534 2748
rect 10590 2746 10614 2748
rect 10670 2746 10676 2748
rect 10430 2694 10432 2746
rect 10612 2694 10614 2746
rect 10368 2692 10374 2694
rect 10430 2692 10454 2694
rect 10510 2692 10534 2694
rect 10590 2692 10614 2694
rect 10670 2692 10676 2694
rect 10368 2683 10676 2692
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 5646 2204 5954 2213
rect 5646 2202 5652 2204
rect 5708 2202 5732 2204
rect 5788 2202 5812 2204
rect 5868 2202 5892 2204
rect 5948 2202 5954 2204
rect 5708 2150 5710 2202
rect 5890 2150 5892 2202
rect 5646 2148 5652 2150
rect 5708 2148 5732 2150
rect 5788 2148 5812 2150
rect 5868 2148 5892 2150
rect 5948 2148 5954 2150
rect 5646 2139 5954 2148
rect 8337 2204 8645 2213
rect 8337 2202 8343 2204
rect 8399 2202 8423 2204
rect 8479 2202 8503 2204
rect 8559 2202 8583 2204
rect 8639 2202 8645 2204
rect 8399 2150 8401 2202
rect 8581 2150 8583 2202
rect 8337 2148 8343 2150
rect 8399 2148 8423 2150
rect 8479 2148 8503 2150
rect 8559 2148 8583 2150
rect 8639 2148 8645 2150
rect 8337 2139 8645 2148
rect 8404 870 8524 898
rect 8404 800 8432 870
rect 5276 734 5488 762
rect 8390 0 8446 800
rect 8496 762 8524 870
rect 8772 762 8800 2246
rect 10704 1494 10732 2790
rect 10796 2446 10824 7686
rect 11028 7644 11336 7653
rect 11028 7642 11034 7644
rect 11090 7642 11114 7644
rect 11170 7642 11194 7644
rect 11250 7642 11274 7644
rect 11330 7642 11336 7644
rect 11090 7590 11092 7642
rect 11272 7590 11274 7642
rect 11028 7588 11034 7590
rect 11090 7588 11114 7590
rect 11170 7588 11194 7590
rect 11250 7588 11274 7590
rect 11330 7588 11336 7590
rect 11028 7579 11336 7588
rect 11028 6556 11336 6565
rect 11028 6554 11034 6556
rect 11090 6554 11114 6556
rect 11170 6554 11194 6556
rect 11250 6554 11274 6556
rect 11330 6554 11336 6556
rect 11090 6502 11092 6554
rect 11272 6502 11274 6554
rect 11028 6500 11034 6502
rect 11090 6500 11114 6502
rect 11170 6500 11194 6502
rect 11250 6500 11274 6502
rect 11330 6500 11336 6502
rect 11028 6491 11336 6500
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10888 5914 10916 6258
rect 11794 6216 11850 6225
rect 11794 6151 11850 6160
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 11808 5710 11836 6151
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11028 5468 11336 5477
rect 11028 5466 11034 5468
rect 11090 5466 11114 5468
rect 11170 5466 11194 5468
rect 11250 5466 11274 5468
rect 11330 5466 11336 5468
rect 11090 5414 11092 5466
rect 11272 5414 11274 5466
rect 11028 5412 11034 5414
rect 11090 5412 11114 5414
rect 11170 5412 11194 5414
rect 11250 5412 11274 5414
rect 11330 5412 11336 5414
rect 11028 5403 11336 5412
rect 11028 4380 11336 4389
rect 11028 4378 11034 4380
rect 11090 4378 11114 4380
rect 11170 4378 11194 4380
rect 11250 4378 11274 4380
rect 11330 4378 11336 4380
rect 11090 4326 11092 4378
rect 11272 4326 11274 4378
rect 11028 4324 11034 4326
rect 11090 4324 11114 4326
rect 11170 4324 11194 4326
rect 11250 4324 11274 4326
rect 11330 4324 11336 4326
rect 11028 4315 11336 4324
rect 11028 3292 11336 3301
rect 11028 3290 11034 3292
rect 11090 3290 11114 3292
rect 11170 3290 11194 3292
rect 11250 3290 11274 3292
rect 11330 3290 11336 3292
rect 11090 3238 11092 3290
rect 11272 3238 11274 3290
rect 11028 3236 11034 3238
rect 11090 3236 11114 3238
rect 11170 3236 11194 3238
rect 11250 3236 11274 3238
rect 11330 3236 11336 3238
rect 11028 3227 11336 3236
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10692 1488 10744 1494
rect 10692 1430 10744 1436
rect 10888 785 10916 2246
rect 11028 2204 11336 2213
rect 11028 2202 11034 2204
rect 11090 2202 11114 2204
rect 11170 2202 11194 2204
rect 11250 2202 11274 2204
rect 11330 2202 11336 2204
rect 11090 2150 11092 2202
rect 11272 2150 11274 2202
rect 11028 2148 11034 2150
rect 11090 2148 11114 2150
rect 11170 2148 11194 2150
rect 11250 2148 11274 2150
rect 11330 2148 11336 2150
rect 11028 2139 11336 2148
rect 10968 1488 11020 1494
rect 10968 1430 11020 1436
rect 10980 800 11008 1430
rect 8496 734 8800 762
rect 10874 776 10930 785
rect 10874 711 10930 720
rect 10966 0 11022 800
<< via2 >>
rect 1398 14048 1454 14104
rect 2301 12538 2357 12540
rect 2381 12538 2437 12540
rect 2461 12538 2517 12540
rect 2541 12538 2597 12540
rect 2301 12486 2347 12538
rect 2347 12486 2357 12538
rect 2381 12486 2411 12538
rect 2411 12486 2423 12538
rect 2423 12486 2437 12538
rect 2461 12486 2475 12538
rect 2475 12486 2487 12538
rect 2487 12486 2517 12538
rect 2541 12486 2551 12538
rect 2551 12486 2597 12538
rect 2301 12484 2357 12486
rect 2381 12484 2437 12486
rect 2461 12484 2517 12486
rect 2541 12484 2597 12486
rect 4992 12538 5048 12540
rect 5072 12538 5128 12540
rect 5152 12538 5208 12540
rect 5232 12538 5288 12540
rect 4992 12486 5038 12538
rect 5038 12486 5048 12538
rect 5072 12486 5102 12538
rect 5102 12486 5114 12538
rect 5114 12486 5128 12538
rect 5152 12486 5166 12538
rect 5166 12486 5178 12538
rect 5178 12486 5208 12538
rect 5232 12486 5242 12538
rect 5242 12486 5288 12538
rect 4992 12484 5048 12486
rect 5072 12484 5128 12486
rect 5152 12484 5208 12486
rect 5232 12484 5288 12486
rect 7683 12538 7739 12540
rect 7763 12538 7819 12540
rect 7843 12538 7899 12540
rect 7923 12538 7979 12540
rect 7683 12486 7729 12538
rect 7729 12486 7739 12538
rect 7763 12486 7793 12538
rect 7793 12486 7805 12538
rect 7805 12486 7819 12538
rect 7843 12486 7857 12538
rect 7857 12486 7869 12538
rect 7869 12486 7899 12538
rect 7923 12486 7933 12538
rect 7933 12486 7979 12538
rect 7683 12484 7739 12486
rect 7763 12484 7819 12486
rect 7843 12484 7899 12486
rect 7923 12484 7979 12486
rect 10374 12538 10430 12540
rect 10454 12538 10510 12540
rect 10534 12538 10590 12540
rect 10614 12538 10670 12540
rect 10374 12486 10420 12538
rect 10420 12486 10430 12538
rect 10454 12486 10484 12538
rect 10484 12486 10496 12538
rect 10496 12486 10510 12538
rect 10534 12486 10548 12538
rect 10548 12486 10560 12538
rect 10560 12486 10590 12538
rect 10614 12486 10624 12538
rect 10624 12486 10670 12538
rect 10374 12484 10430 12486
rect 10454 12484 10510 12486
rect 10534 12484 10590 12486
rect 10614 12484 10670 12486
rect 11242 12280 11298 12336
rect 938 11600 994 11656
rect 2961 11994 3017 11996
rect 3041 11994 3097 11996
rect 3121 11994 3177 11996
rect 3201 11994 3257 11996
rect 2961 11942 3007 11994
rect 3007 11942 3017 11994
rect 3041 11942 3071 11994
rect 3071 11942 3083 11994
rect 3083 11942 3097 11994
rect 3121 11942 3135 11994
rect 3135 11942 3147 11994
rect 3147 11942 3177 11994
rect 3201 11942 3211 11994
rect 3211 11942 3257 11994
rect 2961 11940 3017 11942
rect 3041 11940 3097 11942
rect 3121 11940 3177 11942
rect 3201 11940 3257 11942
rect 2301 11450 2357 11452
rect 2381 11450 2437 11452
rect 2461 11450 2517 11452
rect 2541 11450 2597 11452
rect 2301 11398 2347 11450
rect 2347 11398 2357 11450
rect 2381 11398 2411 11450
rect 2411 11398 2423 11450
rect 2423 11398 2437 11450
rect 2461 11398 2475 11450
rect 2475 11398 2487 11450
rect 2487 11398 2517 11450
rect 2541 11398 2551 11450
rect 2551 11398 2597 11450
rect 2301 11396 2357 11398
rect 2381 11396 2437 11398
rect 2461 11396 2517 11398
rect 2541 11396 2597 11398
rect 2502 10668 2558 10704
rect 2502 10648 2504 10668
rect 2504 10648 2556 10668
rect 2556 10648 2558 10668
rect 2961 10906 3017 10908
rect 3041 10906 3097 10908
rect 3121 10906 3177 10908
rect 3201 10906 3257 10908
rect 2961 10854 3007 10906
rect 3007 10854 3017 10906
rect 3041 10854 3071 10906
rect 3071 10854 3083 10906
rect 3083 10854 3097 10906
rect 3121 10854 3135 10906
rect 3135 10854 3147 10906
rect 3147 10854 3177 10906
rect 3201 10854 3211 10906
rect 3211 10854 3257 10906
rect 2961 10852 3017 10854
rect 3041 10852 3097 10854
rect 3121 10852 3177 10854
rect 3201 10852 3257 10854
rect 2301 10362 2357 10364
rect 2381 10362 2437 10364
rect 2461 10362 2517 10364
rect 2541 10362 2597 10364
rect 2301 10310 2347 10362
rect 2347 10310 2357 10362
rect 2381 10310 2411 10362
rect 2411 10310 2423 10362
rect 2423 10310 2437 10362
rect 2461 10310 2475 10362
rect 2475 10310 2487 10362
rect 2487 10310 2517 10362
rect 2541 10310 2551 10362
rect 2551 10310 2597 10362
rect 2301 10308 2357 10310
rect 2381 10308 2437 10310
rect 2461 10308 2517 10310
rect 2541 10308 2597 10310
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 2961 9818 3017 9820
rect 3041 9818 3097 9820
rect 3121 9818 3177 9820
rect 3201 9818 3257 9820
rect 2961 9766 3007 9818
rect 3007 9766 3017 9818
rect 3041 9766 3071 9818
rect 3071 9766 3083 9818
rect 3083 9766 3097 9818
rect 3121 9766 3135 9818
rect 3135 9766 3147 9818
rect 3147 9766 3177 9818
rect 3201 9766 3211 9818
rect 3211 9766 3257 9818
rect 2961 9764 3017 9766
rect 3041 9764 3097 9766
rect 3121 9764 3177 9766
rect 3201 9764 3257 9766
rect 2301 9274 2357 9276
rect 2381 9274 2437 9276
rect 2461 9274 2517 9276
rect 2541 9274 2597 9276
rect 2301 9222 2347 9274
rect 2347 9222 2357 9274
rect 2381 9222 2411 9274
rect 2411 9222 2423 9274
rect 2423 9222 2437 9274
rect 2461 9222 2475 9274
rect 2475 9222 2487 9274
rect 2487 9222 2517 9274
rect 2541 9222 2551 9274
rect 2551 9222 2597 9274
rect 2301 9220 2357 9222
rect 2381 9220 2437 9222
rect 2461 9220 2517 9222
rect 2541 9220 2597 9222
rect 938 5480 994 5536
rect 938 2760 994 2816
rect 5652 11994 5708 11996
rect 5732 11994 5788 11996
rect 5812 11994 5868 11996
rect 5892 11994 5948 11996
rect 5652 11942 5698 11994
rect 5698 11942 5708 11994
rect 5732 11942 5762 11994
rect 5762 11942 5774 11994
rect 5774 11942 5788 11994
rect 5812 11942 5826 11994
rect 5826 11942 5838 11994
rect 5838 11942 5868 11994
rect 5892 11942 5902 11994
rect 5902 11942 5948 11994
rect 5652 11940 5708 11942
rect 5732 11940 5788 11942
rect 5812 11940 5868 11942
rect 5892 11940 5948 11942
rect 2961 8730 3017 8732
rect 3041 8730 3097 8732
rect 3121 8730 3177 8732
rect 3201 8730 3257 8732
rect 2961 8678 3007 8730
rect 3007 8678 3017 8730
rect 3041 8678 3071 8730
rect 3071 8678 3083 8730
rect 3083 8678 3097 8730
rect 3121 8678 3135 8730
rect 3135 8678 3147 8730
rect 3147 8678 3177 8730
rect 3201 8678 3211 8730
rect 3211 8678 3257 8730
rect 2961 8676 3017 8678
rect 3041 8676 3097 8678
rect 3121 8676 3177 8678
rect 3201 8676 3257 8678
rect 2301 8186 2357 8188
rect 2381 8186 2437 8188
rect 2461 8186 2517 8188
rect 2541 8186 2597 8188
rect 2301 8134 2347 8186
rect 2347 8134 2357 8186
rect 2381 8134 2411 8186
rect 2411 8134 2423 8186
rect 2423 8134 2437 8186
rect 2461 8134 2475 8186
rect 2475 8134 2487 8186
rect 2487 8134 2517 8186
rect 2541 8134 2551 8186
rect 2551 8134 2597 8186
rect 2301 8132 2357 8134
rect 2381 8132 2437 8134
rect 2461 8132 2517 8134
rect 2541 8132 2597 8134
rect 4992 11450 5048 11452
rect 5072 11450 5128 11452
rect 5152 11450 5208 11452
rect 5232 11450 5288 11452
rect 4992 11398 5038 11450
rect 5038 11398 5048 11450
rect 5072 11398 5102 11450
rect 5102 11398 5114 11450
rect 5114 11398 5128 11450
rect 5152 11398 5166 11450
rect 5166 11398 5178 11450
rect 5178 11398 5208 11450
rect 5232 11398 5242 11450
rect 5242 11398 5288 11450
rect 4992 11396 5048 11398
rect 5072 11396 5128 11398
rect 5152 11396 5208 11398
rect 5232 11396 5288 11398
rect 5446 10648 5502 10704
rect 4992 10362 5048 10364
rect 5072 10362 5128 10364
rect 5152 10362 5208 10364
rect 5232 10362 5288 10364
rect 4992 10310 5038 10362
rect 5038 10310 5048 10362
rect 5072 10310 5102 10362
rect 5102 10310 5114 10362
rect 5114 10310 5128 10362
rect 5152 10310 5166 10362
rect 5166 10310 5178 10362
rect 5178 10310 5208 10362
rect 5232 10310 5242 10362
rect 5242 10310 5288 10362
rect 4992 10308 5048 10310
rect 5072 10308 5128 10310
rect 5152 10308 5208 10310
rect 5232 10308 5288 10310
rect 7683 11450 7739 11452
rect 7763 11450 7819 11452
rect 7843 11450 7899 11452
rect 7923 11450 7979 11452
rect 7683 11398 7729 11450
rect 7729 11398 7739 11450
rect 7763 11398 7793 11450
rect 7793 11398 7805 11450
rect 7805 11398 7819 11450
rect 7843 11398 7857 11450
rect 7857 11398 7869 11450
rect 7869 11398 7899 11450
rect 7923 11398 7933 11450
rect 7933 11398 7979 11450
rect 7683 11396 7739 11398
rect 7763 11396 7819 11398
rect 7843 11396 7899 11398
rect 7923 11396 7979 11398
rect 5652 10906 5708 10908
rect 5732 10906 5788 10908
rect 5812 10906 5868 10908
rect 5892 10906 5948 10908
rect 5652 10854 5698 10906
rect 5698 10854 5708 10906
rect 5732 10854 5762 10906
rect 5762 10854 5774 10906
rect 5774 10854 5788 10906
rect 5812 10854 5826 10906
rect 5826 10854 5838 10906
rect 5838 10854 5868 10906
rect 5892 10854 5902 10906
rect 5902 10854 5948 10906
rect 5652 10852 5708 10854
rect 5732 10852 5788 10854
rect 5812 10852 5868 10854
rect 5892 10852 5948 10854
rect 2961 7642 3017 7644
rect 3041 7642 3097 7644
rect 3121 7642 3177 7644
rect 3201 7642 3257 7644
rect 2961 7590 3007 7642
rect 3007 7590 3017 7642
rect 3041 7590 3071 7642
rect 3071 7590 3083 7642
rect 3083 7590 3097 7642
rect 3121 7590 3135 7642
rect 3135 7590 3147 7642
rect 3147 7590 3177 7642
rect 3201 7590 3211 7642
rect 3211 7590 3257 7642
rect 2961 7588 3017 7590
rect 3041 7588 3097 7590
rect 3121 7588 3177 7590
rect 3201 7588 3257 7590
rect 2301 7098 2357 7100
rect 2381 7098 2437 7100
rect 2461 7098 2517 7100
rect 2541 7098 2597 7100
rect 2301 7046 2347 7098
rect 2347 7046 2357 7098
rect 2381 7046 2411 7098
rect 2411 7046 2423 7098
rect 2423 7046 2437 7098
rect 2461 7046 2475 7098
rect 2475 7046 2487 7098
rect 2487 7046 2517 7098
rect 2541 7046 2551 7098
rect 2551 7046 2597 7098
rect 2301 7044 2357 7046
rect 2381 7044 2437 7046
rect 2461 7044 2517 7046
rect 2541 7044 2597 7046
rect 2961 6554 3017 6556
rect 3041 6554 3097 6556
rect 3121 6554 3177 6556
rect 3201 6554 3257 6556
rect 2961 6502 3007 6554
rect 3007 6502 3017 6554
rect 3041 6502 3071 6554
rect 3071 6502 3083 6554
rect 3083 6502 3097 6554
rect 3121 6502 3135 6554
rect 3135 6502 3147 6554
rect 3147 6502 3177 6554
rect 3201 6502 3211 6554
rect 3211 6502 3257 6554
rect 2961 6500 3017 6502
rect 3041 6500 3097 6502
rect 3121 6500 3177 6502
rect 3201 6500 3257 6502
rect 2301 6010 2357 6012
rect 2381 6010 2437 6012
rect 2461 6010 2517 6012
rect 2541 6010 2597 6012
rect 2301 5958 2347 6010
rect 2347 5958 2357 6010
rect 2381 5958 2411 6010
rect 2411 5958 2423 6010
rect 2423 5958 2437 6010
rect 2461 5958 2475 6010
rect 2475 5958 2487 6010
rect 2487 5958 2517 6010
rect 2541 5958 2551 6010
rect 2551 5958 2597 6010
rect 2301 5956 2357 5958
rect 2381 5956 2437 5958
rect 2461 5956 2517 5958
rect 2541 5956 2597 5958
rect 2961 5466 3017 5468
rect 3041 5466 3097 5468
rect 3121 5466 3177 5468
rect 3201 5466 3257 5468
rect 2961 5414 3007 5466
rect 3007 5414 3017 5466
rect 3041 5414 3071 5466
rect 3071 5414 3083 5466
rect 3083 5414 3097 5466
rect 3121 5414 3135 5466
rect 3135 5414 3147 5466
rect 3147 5414 3177 5466
rect 3201 5414 3211 5466
rect 3211 5414 3257 5466
rect 2961 5412 3017 5414
rect 3041 5412 3097 5414
rect 3121 5412 3177 5414
rect 3201 5412 3257 5414
rect 2301 4922 2357 4924
rect 2381 4922 2437 4924
rect 2461 4922 2517 4924
rect 2541 4922 2597 4924
rect 2301 4870 2347 4922
rect 2347 4870 2357 4922
rect 2381 4870 2411 4922
rect 2411 4870 2423 4922
rect 2423 4870 2437 4922
rect 2461 4870 2475 4922
rect 2475 4870 2487 4922
rect 2487 4870 2517 4922
rect 2541 4870 2551 4922
rect 2551 4870 2597 4922
rect 2301 4868 2357 4870
rect 2381 4868 2437 4870
rect 2461 4868 2517 4870
rect 2541 4868 2597 4870
rect 2301 3834 2357 3836
rect 2381 3834 2437 3836
rect 2461 3834 2517 3836
rect 2541 3834 2597 3836
rect 2301 3782 2347 3834
rect 2347 3782 2357 3834
rect 2381 3782 2411 3834
rect 2411 3782 2423 3834
rect 2423 3782 2437 3834
rect 2461 3782 2475 3834
rect 2475 3782 2487 3834
rect 2487 3782 2517 3834
rect 2541 3782 2551 3834
rect 2551 3782 2597 3834
rect 2301 3780 2357 3782
rect 2381 3780 2437 3782
rect 2461 3780 2517 3782
rect 2541 3780 2597 3782
rect 2961 4378 3017 4380
rect 3041 4378 3097 4380
rect 3121 4378 3177 4380
rect 3201 4378 3257 4380
rect 2961 4326 3007 4378
rect 3007 4326 3017 4378
rect 3041 4326 3071 4378
rect 3071 4326 3083 4378
rect 3083 4326 3097 4378
rect 3121 4326 3135 4378
rect 3135 4326 3147 4378
rect 3147 4326 3177 4378
rect 3201 4326 3211 4378
rect 3211 4326 3257 4378
rect 2961 4324 3017 4326
rect 3041 4324 3097 4326
rect 3121 4324 3177 4326
rect 3201 4324 3257 4326
rect 2961 3290 3017 3292
rect 3041 3290 3097 3292
rect 3121 3290 3177 3292
rect 3201 3290 3257 3292
rect 2961 3238 3007 3290
rect 3007 3238 3017 3290
rect 3041 3238 3071 3290
rect 3071 3238 3083 3290
rect 3083 3238 3097 3290
rect 3121 3238 3135 3290
rect 3135 3238 3147 3290
rect 3147 3238 3177 3290
rect 3201 3238 3211 3290
rect 3211 3238 3257 3290
rect 2961 3236 3017 3238
rect 3041 3236 3097 3238
rect 3121 3236 3177 3238
rect 3201 3236 3257 3238
rect 2301 2746 2357 2748
rect 2381 2746 2437 2748
rect 2461 2746 2517 2748
rect 2541 2746 2597 2748
rect 2301 2694 2347 2746
rect 2347 2694 2357 2746
rect 2381 2694 2411 2746
rect 2411 2694 2423 2746
rect 2423 2694 2437 2746
rect 2461 2694 2475 2746
rect 2475 2694 2487 2746
rect 2487 2694 2517 2746
rect 2541 2694 2551 2746
rect 2551 2694 2597 2746
rect 2301 2692 2357 2694
rect 2381 2692 2437 2694
rect 2461 2692 2517 2694
rect 2541 2692 2597 2694
rect 7683 10362 7739 10364
rect 7763 10362 7819 10364
rect 7843 10362 7899 10364
rect 7923 10362 7979 10364
rect 7683 10310 7729 10362
rect 7729 10310 7739 10362
rect 7763 10310 7793 10362
rect 7793 10310 7805 10362
rect 7805 10310 7819 10362
rect 7843 10310 7857 10362
rect 7857 10310 7869 10362
rect 7869 10310 7899 10362
rect 7923 10310 7933 10362
rect 7933 10310 7979 10362
rect 7683 10308 7739 10310
rect 7763 10308 7819 10310
rect 7843 10308 7899 10310
rect 7923 10308 7979 10310
rect 5652 9818 5708 9820
rect 5732 9818 5788 9820
rect 5812 9818 5868 9820
rect 5892 9818 5948 9820
rect 5652 9766 5698 9818
rect 5698 9766 5708 9818
rect 5732 9766 5762 9818
rect 5762 9766 5774 9818
rect 5774 9766 5788 9818
rect 5812 9766 5826 9818
rect 5826 9766 5838 9818
rect 5838 9766 5868 9818
rect 5892 9766 5902 9818
rect 5902 9766 5948 9818
rect 5652 9764 5708 9766
rect 5732 9764 5788 9766
rect 5812 9764 5868 9766
rect 5892 9764 5948 9766
rect 4992 9274 5048 9276
rect 5072 9274 5128 9276
rect 5152 9274 5208 9276
rect 5232 9274 5288 9276
rect 4992 9222 5038 9274
rect 5038 9222 5048 9274
rect 5072 9222 5102 9274
rect 5102 9222 5114 9274
rect 5114 9222 5128 9274
rect 5152 9222 5166 9274
rect 5166 9222 5178 9274
rect 5178 9222 5208 9274
rect 5232 9222 5242 9274
rect 5242 9222 5288 9274
rect 4992 9220 5048 9222
rect 5072 9220 5128 9222
rect 5152 9220 5208 9222
rect 5232 9220 5288 9222
rect 4992 8186 5048 8188
rect 5072 8186 5128 8188
rect 5152 8186 5208 8188
rect 5232 8186 5288 8188
rect 4992 8134 5038 8186
rect 5038 8134 5048 8186
rect 5072 8134 5102 8186
rect 5102 8134 5114 8186
rect 5114 8134 5128 8186
rect 5152 8134 5166 8186
rect 5166 8134 5178 8186
rect 5178 8134 5208 8186
rect 5232 8134 5242 8186
rect 5242 8134 5288 8186
rect 4992 8132 5048 8134
rect 5072 8132 5128 8134
rect 5152 8132 5208 8134
rect 5232 8132 5288 8134
rect 4992 7098 5048 7100
rect 5072 7098 5128 7100
rect 5152 7098 5208 7100
rect 5232 7098 5288 7100
rect 4992 7046 5038 7098
rect 5038 7046 5048 7098
rect 5072 7046 5102 7098
rect 5102 7046 5114 7098
rect 5114 7046 5128 7098
rect 5152 7046 5166 7098
rect 5166 7046 5178 7098
rect 5178 7046 5208 7098
rect 5232 7046 5242 7098
rect 5242 7046 5288 7098
rect 4992 7044 5048 7046
rect 5072 7044 5128 7046
rect 5152 7044 5208 7046
rect 5232 7044 5288 7046
rect 7683 9274 7739 9276
rect 7763 9274 7819 9276
rect 7843 9274 7899 9276
rect 7923 9274 7979 9276
rect 7683 9222 7729 9274
rect 7729 9222 7739 9274
rect 7763 9222 7793 9274
rect 7793 9222 7805 9274
rect 7805 9222 7819 9274
rect 7843 9222 7857 9274
rect 7857 9222 7869 9274
rect 7869 9222 7899 9274
rect 7923 9222 7933 9274
rect 7933 9222 7979 9274
rect 7683 9220 7739 9222
rect 7763 9220 7819 9222
rect 7843 9220 7899 9222
rect 7923 9220 7979 9222
rect 5652 8730 5708 8732
rect 5732 8730 5788 8732
rect 5812 8730 5868 8732
rect 5892 8730 5948 8732
rect 5652 8678 5698 8730
rect 5698 8678 5708 8730
rect 5732 8678 5762 8730
rect 5762 8678 5774 8730
rect 5774 8678 5788 8730
rect 5812 8678 5826 8730
rect 5826 8678 5838 8730
rect 5838 8678 5868 8730
rect 5892 8678 5902 8730
rect 5902 8678 5948 8730
rect 5652 8676 5708 8678
rect 5732 8676 5788 8678
rect 5812 8676 5868 8678
rect 5892 8676 5948 8678
rect 5652 7642 5708 7644
rect 5732 7642 5788 7644
rect 5812 7642 5868 7644
rect 5892 7642 5948 7644
rect 5652 7590 5698 7642
rect 5698 7590 5708 7642
rect 5732 7590 5762 7642
rect 5762 7590 5774 7642
rect 5774 7590 5788 7642
rect 5812 7590 5826 7642
rect 5826 7590 5838 7642
rect 5838 7590 5868 7642
rect 5892 7590 5902 7642
rect 5902 7590 5948 7642
rect 5652 7588 5708 7590
rect 5732 7588 5788 7590
rect 5812 7588 5868 7590
rect 5892 7588 5948 7590
rect 5652 6554 5708 6556
rect 5732 6554 5788 6556
rect 5812 6554 5868 6556
rect 5892 6554 5948 6556
rect 5652 6502 5698 6554
rect 5698 6502 5708 6554
rect 5732 6502 5762 6554
rect 5762 6502 5774 6554
rect 5774 6502 5788 6554
rect 5812 6502 5826 6554
rect 5826 6502 5838 6554
rect 5838 6502 5868 6554
rect 5892 6502 5902 6554
rect 5902 6502 5948 6554
rect 5652 6500 5708 6502
rect 5732 6500 5788 6502
rect 5812 6500 5868 6502
rect 5892 6500 5948 6502
rect 4992 6010 5048 6012
rect 5072 6010 5128 6012
rect 5152 6010 5208 6012
rect 5232 6010 5288 6012
rect 4992 5958 5038 6010
rect 5038 5958 5048 6010
rect 5072 5958 5102 6010
rect 5102 5958 5114 6010
rect 5114 5958 5128 6010
rect 5152 5958 5166 6010
rect 5166 5958 5178 6010
rect 5178 5958 5208 6010
rect 5232 5958 5242 6010
rect 5242 5958 5288 6010
rect 4992 5956 5048 5958
rect 5072 5956 5128 5958
rect 5152 5956 5208 5958
rect 5232 5956 5288 5958
rect 4992 4922 5048 4924
rect 5072 4922 5128 4924
rect 5152 4922 5208 4924
rect 5232 4922 5288 4924
rect 4992 4870 5038 4922
rect 5038 4870 5048 4922
rect 5072 4870 5102 4922
rect 5102 4870 5114 4922
rect 5114 4870 5128 4922
rect 5152 4870 5166 4922
rect 5166 4870 5178 4922
rect 5178 4870 5208 4922
rect 5232 4870 5242 4922
rect 5242 4870 5288 4922
rect 4992 4868 5048 4870
rect 5072 4868 5128 4870
rect 5152 4868 5208 4870
rect 5232 4868 5288 4870
rect 5652 5466 5708 5468
rect 5732 5466 5788 5468
rect 5812 5466 5868 5468
rect 5892 5466 5948 5468
rect 5652 5414 5698 5466
rect 5698 5414 5708 5466
rect 5732 5414 5762 5466
rect 5762 5414 5774 5466
rect 5774 5414 5788 5466
rect 5812 5414 5826 5466
rect 5826 5414 5838 5466
rect 5838 5414 5868 5466
rect 5892 5414 5902 5466
rect 5902 5414 5948 5466
rect 5652 5412 5708 5414
rect 5732 5412 5788 5414
rect 5812 5412 5868 5414
rect 5892 5412 5948 5414
rect 5652 4378 5708 4380
rect 5732 4378 5788 4380
rect 5812 4378 5868 4380
rect 5892 4378 5948 4380
rect 5652 4326 5698 4378
rect 5698 4326 5708 4378
rect 5732 4326 5762 4378
rect 5762 4326 5774 4378
rect 5774 4326 5788 4378
rect 5812 4326 5826 4378
rect 5826 4326 5838 4378
rect 5838 4326 5868 4378
rect 5892 4326 5902 4378
rect 5902 4326 5948 4378
rect 5652 4324 5708 4326
rect 5732 4324 5788 4326
rect 5812 4324 5868 4326
rect 5892 4324 5948 4326
rect 6274 6704 6330 6760
rect 7683 8186 7739 8188
rect 7763 8186 7819 8188
rect 7843 8186 7899 8188
rect 7923 8186 7979 8188
rect 7683 8134 7729 8186
rect 7729 8134 7739 8186
rect 7763 8134 7793 8186
rect 7793 8134 7805 8186
rect 7805 8134 7819 8186
rect 7843 8134 7857 8186
rect 7857 8134 7869 8186
rect 7869 8134 7899 8186
rect 7923 8134 7933 8186
rect 7933 8134 7979 8186
rect 7683 8132 7739 8134
rect 7763 8132 7819 8134
rect 7843 8132 7899 8134
rect 7923 8132 7979 8134
rect 6918 6976 6974 7032
rect 7683 7098 7739 7100
rect 7763 7098 7819 7100
rect 7843 7098 7899 7100
rect 7923 7098 7979 7100
rect 7683 7046 7729 7098
rect 7729 7046 7739 7098
rect 7763 7046 7793 7098
rect 7793 7046 7805 7098
rect 7805 7046 7819 7098
rect 7843 7046 7857 7098
rect 7857 7046 7869 7098
rect 7869 7046 7899 7098
rect 7923 7046 7933 7098
rect 7933 7046 7979 7098
rect 7683 7044 7739 7046
rect 7763 7044 7819 7046
rect 7843 7044 7899 7046
rect 7923 7044 7979 7046
rect 6918 6296 6974 6352
rect 7562 6704 7618 6760
rect 8343 11994 8399 11996
rect 8423 11994 8479 11996
rect 8503 11994 8559 11996
rect 8583 11994 8639 11996
rect 8343 11942 8389 11994
rect 8389 11942 8399 11994
rect 8423 11942 8453 11994
rect 8453 11942 8465 11994
rect 8465 11942 8479 11994
rect 8503 11942 8517 11994
rect 8517 11942 8529 11994
rect 8529 11942 8559 11994
rect 8583 11942 8593 11994
rect 8593 11942 8639 11994
rect 8343 11940 8399 11942
rect 8423 11940 8479 11942
rect 8503 11940 8559 11942
rect 8583 11940 8639 11942
rect 11034 11994 11090 11996
rect 11114 11994 11170 11996
rect 11194 11994 11250 11996
rect 11274 11994 11330 11996
rect 11034 11942 11080 11994
rect 11080 11942 11090 11994
rect 11114 11942 11144 11994
rect 11144 11942 11156 11994
rect 11156 11942 11170 11994
rect 11194 11942 11208 11994
rect 11208 11942 11220 11994
rect 11220 11942 11250 11994
rect 11274 11942 11284 11994
rect 11284 11942 11330 11994
rect 11034 11940 11090 11942
rect 11114 11940 11170 11942
rect 11194 11940 11250 11942
rect 11274 11940 11330 11942
rect 8343 10906 8399 10908
rect 8423 10906 8479 10908
rect 8503 10906 8559 10908
rect 8583 10906 8639 10908
rect 8343 10854 8389 10906
rect 8389 10854 8399 10906
rect 8423 10854 8453 10906
rect 8453 10854 8465 10906
rect 8465 10854 8479 10906
rect 8503 10854 8517 10906
rect 8517 10854 8529 10906
rect 8529 10854 8559 10906
rect 8583 10854 8593 10906
rect 8593 10854 8639 10906
rect 8343 10852 8399 10854
rect 8423 10852 8479 10854
rect 8503 10852 8559 10854
rect 8583 10852 8639 10854
rect 10374 11450 10430 11452
rect 10454 11450 10510 11452
rect 10534 11450 10590 11452
rect 10614 11450 10670 11452
rect 10374 11398 10420 11450
rect 10420 11398 10430 11450
rect 10454 11398 10484 11450
rect 10484 11398 10496 11450
rect 10496 11398 10510 11450
rect 10534 11398 10548 11450
rect 10548 11398 10560 11450
rect 10560 11398 10590 11450
rect 10614 11398 10624 11450
rect 10624 11398 10670 11450
rect 10374 11396 10430 11398
rect 10454 11396 10510 11398
rect 10534 11396 10590 11398
rect 10614 11396 10670 11398
rect 8343 9818 8399 9820
rect 8423 9818 8479 9820
rect 8503 9818 8559 9820
rect 8583 9818 8639 9820
rect 8343 9766 8389 9818
rect 8389 9766 8399 9818
rect 8423 9766 8453 9818
rect 8453 9766 8465 9818
rect 8465 9766 8479 9818
rect 8503 9766 8517 9818
rect 8517 9766 8529 9818
rect 8529 9766 8559 9818
rect 8583 9766 8593 9818
rect 8593 9766 8639 9818
rect 8343 9764 8399 9766
rect 8423 9764 8479 9766
rect 8503 9764 8559 9766
rect 8583 9764 8639 9766
rect 8343 8730 8399 8732
rect 8423 8730 8479 8732
rect 8503 8730 8559 8732
rect 8583 8730 8639 8732
rect 8343 8678 8389 8730
rect 8389 8678 8399 8730
rect 8423 8678 8453 8730
rect 8453 8678 8465 8730
rect 8465 8678 8479 8730
rect 8503 8678 8517 8730
rect 8517 8678 8529 8730
rect 8529 8678 8559 8730
rect 8583 8678 8593 8730
rect 8593 8678 8639 8730
rect 8343 8676 8399 8678
rect 8423 8676 8479 8678
rect 8503 8676 8559 8678
rect 8583 8676 8639 8678
rect 8343 7642 8399 7644
rect 8423 7642 8479 7644
rect 8503 7642 8559 7644
rect 8583 7642 8639 7644
rect 8343 7590 8389 7642
rect 8389 7590 8399 7642
rect 8423 7590 8453 7642
rect 8453 7590 8465 7642
rect 8465 7590 8479 7642
rect 8503 7590 8517 7642
rect 8517 7590 8529 7642
rect 8529 7590 8559 7642
rect 8583 7590 8593 7642
rect 8593 7590 8639 7642
rect 8343 7588 8399 7590
rect 8423 7588 8479 7590
rect 8503 7588 8559 7590
rect 8583 7588 8639 7590
rect 8206 6976 8262 7032
rect 8343 6554 8399 6556
rect 8423 6554 8479 6556
rect 8503 6554 8559 6556
rect 8583 6554 8639 6556
rect 8343 6502 8389 6554
rect 8389 6502 8399 6554
rect 8423 6502 8453 6554
rect 8453 6502 8465 6554
rect 8465 6502 8479 6554
rect 8503 6502 8517 6554
rect 8517 6502 8529 6554
rect 8529 6502 8559 6554
rect 8583 6502 8593 6554
rect 8593 6502 8639 6554
rect 8343 6500 8399 6502
rect 8423 6500 8479 6502
rect 8503 6500 8559 6502
rect 8583 6500 8639 6502
rect 7683 6010 7739 6012
rect 7763 6010 7819 6012
rect 7843 6010 7899 6012
rect 7923 6010 7979 6012
rect 7683 5958 7729 6010
rect 7729 5958 7739 6010
rect 7763 5958 7793 6010
rect 7793 5958 7805 6010
rect 7805 5958 7819 6010
rect 7843 5958 7857 6010
rect 7857 5958 7869 6010
rect 7869 5958 7899 6010
rect 7923 5958 7933 6010
rect 7933 5958 7979 6010
rect 7683 5956 7739 5958
rect 7763 5956 7819 5958
rect 7843 5956 7899 5958
rect 7923 5956 7979 5958
rect 6182 3984 6238 4040
rect 4992 3834 5048 3836
rect 5072 3834 5128 3836
rect 5152 3834 5208 3836
rect 5232 3834 5288 3836
rect 4992 3782 5038 3834
rect 5038 3782 5048 3834
rect 5072 3782 5102 3834
rect 5102 3782 5114 3834
rect 5114 3782 5128 3834
rect 5152 3782 5166 3834
rect 5166 3782 5178 3834
rect 5178 3782 5208 3834
rect 5232 3782 5242 3834
rect 5242 3782 5288 3834
rect 4992 3780 5048 3782
rect 5072 3780 5128 3782
rect 5152 3780 5208 3782
rect 5232 3780 5288 3782
rect 5652 3290 5708 3292
rect 5732 3290 5788 3292
rect 5812 3290 5868 3292
rect 5892 3290 5948 3292
rect 5652 3238 5698 3290
rect 5698 3238 5708 3290
rect 5732 3238 5762 3290
rect 5762 3238 5774 3290
rect 5774 3238 5788 3290
rect 5812 3238 5826 3290
rect 5826 3238 5838 3290
rect 5838 3238 5868 3290
rect 5892 3238 5902 3290
rect 5902 3238 5948 3290
rect 5652 3236 5708 3238
rect 5732 3236 5788 3238
rect 5812 3236 5868 3238
rect 5892 3236 5948 3238
rect 4992 2746 5048 2748
rect 5072 2746 5128 2748
rect 5152 2746 5208 2748
rect 5232 2746 5288 2748
rect 4992 2694 5038 2746
rect 5038 2694 5048 2746
rect 5072 2694 5102 2746
rect 5102 2694 5114 2746
rect 5114 2694 5128 2746
rect 5152 2694 5166 2746
rect 5166 2694 5178 2746
rect 5178 2694 5208 2746
rect 5232 2694 5242 2746
rect 5242 2694 5288 2746
rect 4992 2692 5048 2694
rect 5072 2692 5128 2694
rect 5152 2692 5208 2694
rect 5232 2692 5288 2694
rect 2961 2202 3017 2204
rect 3041 2202 3097 2204
rect 3121 2202 3177 2204
rect 3201 2202 3257 2204
rect 2961 2150 3007 2202
rect 3007 2150 3017 2202
rect 3041 2150 3071 2202
rect 3071 2150 3083 2202
rect 3083 2150 3097 2202
rect 3121 2150 3135 2202
rect 3135 2150 3147 2202
rect 3147 2150 3177 2202
rect 3201 2150 3211 2202
rect 3211 2150 3257 2202
rect 2961 2148 3017 2150
rect 3041 2148 3097 2150
rect 3121 2148 3177 2150
rect 3201 2148 3257 2150
rect 7683 4922 7739 4924
rect 7763 4922 7819 4924
rect 7843 4922 7899 4924
rect 7923 4922 7979 4924
rect 7683 4870 7729 4922
rect 7729 4870 7739 4922
rect 7763 4870 7793 4922
rect 7793 4870 7805 4922
rect 7805 4870 7819 4922
rect 7843 4870 7857 4922
rect 7857 4870 7869 4922
rect 7869 4870 7899 4922
rect 7923 4870 7933 4922
rect 7933 4870 7979 4922
rect 7683 4868 7739 4870
rect 7763 4868 7819 4870
rect 7843 4868 7899 4870
rect 7923 4868 7979 4870
rect 7683 3834 7739 3836
rect 7763 3834 7819 3836
rect 7843 3834 7899 3836
rect 7923 3834 7979 3836
rect 7683 3782 7729 3834
rect 7729 3782 7739 3834
rect 7763 3782 7793 3834
rect 7793 3782 7805 3834
rect 7805 3782 7819 3834
rect 7843 3782 7857 3834
rect 7857 3782 7869 3834
rect 7869 3782 7899 3834
rect 7923 3782 7933 3834
rect 7933 3782 7979 3834
rect 7683 3780 7739 3782
rect 7763 3780 7819 3782
rect 7843 3780 7899 3782
rect 7923 3780 7979 3782
rect 8343 5466 8399 5468
rect 8423 5466 8479 5468
rect 8503 5466 8559 5468
rect 8583 5466 8639 5468
rect 8343 5414 8389 5466
rect 8389 5414 8399 5466
rect 8423 5414 8453 5466
rect 8453 5414 8465 5466
rect 8465 5414 8479 5466
rect 8503 5414 8517 5466
rect 8517 5414 8529 5466
rect 8529 5414 8559 5466
rect 8583 5414 8593 5466
rect 8593 5414 8639 5466
rect 8343 5412 8399 5414
rect 8423 5412 8479 5414
rect 8503 5412 8559 5414
rect 8583 5412 8639 5414
rect 9034 6296 9090 6352
rect 11034 10906 11090 10908
rect 11114 10906 11170 10908
rect 11194 10906 11250 10908
rect 11274 10906 11330 10908
rect 11034 10854 11080 10906
rect 11080 10854 11090 10906
rect 11114 10854 11144 10906
rect 11144 10854 11156 10906
rect 11156 10854 11170 10906
rect 11194 10854 11208 10906
rect 11208 10854 11220 10906
rect 11220 10854 11250 10906
rect 11274 10854 11284 10906
rect 11284 10854 11330 10906
rect 11034 10852 11090 10854
rect 11114 10852 11170 10854
rect 11194 10852 11250 10854
rect 11274 10852 11330 10854
rect 10374 10362 10430 10364
rect 10454 10362 10510 10364
rect 10534 10362 10590 10364
rect 10614 10362 10670 10364
rect 10374 10310 10420 10362
rect 10420 10310 10430 10362
rect 10454 10310 10484 10362
rect 10484 10310 10496 10362
rect 10496 10310 10510 10362
rect 10534 10310 10548 10362
rect 10548 10310 10560 10362
rect 10560 10310 10590 10362
rect 10614 10310 10624 10362
rect 10624 10310 10670 10362
rect 10374 10308 10430 10310
rect 10454 10308 10510 10310
rect 10534 10308 10590 10310
rect 10614 10308 10670 10310
rect 10374 9274 10430 9276
rect 10454 9274 10510 9276
rect 10534 9274 10590 9276
rect 10614 9274 10670 9276
rect 10374 9222 10420 9274
rect 10420 9222 10430 9274
rect 10454 9222 10484 9274
rect 10484 9222 10496 9274
rect 10496 9222 10510 9274
rect 10534 9222 10548 9274
rect 10548 9222 10560 9274
rect 10560 9222 10590 9274
rect 10614 9222 10624 9274
rect 10624 9222 10670 9274
rect 10374 9220 10430 9222
rect 10454 9220 10510 9222
rect 10534 9220 10590 9222
rect 10614 9220 10670 9222
rect 10374 8186 10430 8188
rect 10454 8186 10510 8188
rect 10534 8186 10590 8188
rect 10614 8186 10670 8188
rect 10374 8134 10420 8186
rect 10420 8134 10430 8186
rect 10454 8134 10484 8186
rect 10484 8134 10496 8186
rect 10496 8134 10510 8186
rect 10534 8134 10548 8186
rect 10548 8134 10560 8186
rect 10560 8134 10590 8186
rect 10614 8134 10624 8186
rect 10624 8134 10670 8186
rect 10374 8132 10430 8134
rect 10454 8132 10510 8134
rect 10534 8132 10590 8134
rect 10614 8132 10670 8134
rect 11034 9818 11090 9820
rect 11114 9818 11170 9820
rect 11194 9818 11250 9820
rect 11274 9818 11330 9820
rect 11034 9766 11080 9818
rect 11080 9766 11090 9818
rect 11114 9766 11144 9818
rect 11144 9766 11156 9818
rect 11156 9766 11170 9818
rect 11194 9766 11208 9818
rect 11208 9766 11220 9818
rect 11220 9766 11250 9818
rect 11274 9766 11284 9818
rect 11284 9766 11330 9818
rect 11034 9764 11090 9766
rect 11114 9764 11170 9766
rect 11194 9764 11250 9766
rect 11274 9764 11330 9766
rect 12070 9560 12126 9616
rect 11034 8730 11090 8732
rect 11114 8730 11170 8732
rect 11194 8730 11250 8732
rect 11274 8730 11330 8732
rect 11034 8678 11080 8730
rect 11080 8678 11090 8730
rect 11114 8678 11144 8730
rect 11144 8678 11156 8730
rect 11156 8678 11170 8730
rect 11194 8678 11208 8730
rect 11208 8678 11220 8730
rect 11220 8678 11250 8730
rect 11274 8678 11284 8730
rect 11284 8678 11330 8730
rect 11034 8676 11090 8678
rect 11114 8676 11170 8678
rect 11194 8676 11250 8678
rect 11274 8676 11330 8678
rect 10374 7098 10430 7100
rect 10454 7098 10510 7100
rect 10534 7098 10590 7100
rect 10614 7098 10670 7100
rect 10374 7046 10420 7098
rect 10420 7046 10430 7098
rect 10454 7046 10484 7098
rect 10484 7046 10496 7098
rect 10496 7046 10510 7098
rect 10534 7046 10548 7098
rect 10548 7046 10560 7098
rect 10560 7046 10590 7098
rect 10614 7046 10624 7098
rect 10624 7046 10670 7098
rect 10374 7044 10430 7046
rect 10454 7044 10510 7046
rect 10534 7044 10590 7046
rect 10614 7044 10670 7046
rect 8343 4378 8399 4380
rect 8423 4378 8479 4380
rect 8503 4378 8559 4380
rect 8583 4378 8639 4380
rect 8343 4326 8389 4378
rect 8389 4326 8399 4378
rect 8423 4326 8453 4378
rect 8453 4326 8465 4378
rect 8465 4326 8479 4378
rect 8503 4326 8517 4378
rect 8517 4326 8529 4378
rect 8529 4326 8559 4378
rect 8583 4326 8593 4378
rect 8593 4326 8639 4378
rect 8343 4324 8399 4326
rect 8423 4324 8479 4326
rect 8503 4324 8559 4326
rect 8583 4324 8639 4326
rect 7683 2746 7739 2748
rect 7763 2746 7819 2748
rect 7843 2746 7899 2748
rect 7923 2746 7979 2748
rect 7683 2694 7729 2746
rect 7729 2694 7739 2746
rect 7763 2694 7793 2746
rect 7793 2694 7805 2746
rect 7805 2694 7819 2746
rect 7843 2694 7857 2746
rect 7857 2694 7869 2746
rect 7869 2694 7899 2746
rect 7923 2694 7933 2746
rect 7933 2694 7979 2746
rect 7683 2692 7739 2694
rect 7763 2692 7819 2694
rect 7843 2692 7899 2694
rect 7923 2692 7979 2694
rect 8343 3290 8399 3292
rect 8423 3290 8479 3292
rect 8503 3290 8559 3292
rect 8583 3290 8639 3292
rect 8343 3238 8389 3290
rect 8389 3238 8399 3290
rect 8423 3238 8453 3290
rect 8453 3238 8465 3290
rect 8465 3238 8479 3290
rect 8503 3238 8517 3290
rect 8517 3238 8529 3290
rect 8529 3238 8559 3290
rect 8583 3238 8593 3290
rect 8593 3238 8639 3290
rect 8343 3236 8399 3238
rect 8423 3236 8479 3238
rect 8503 3236 8559 3238
rect 8583 3236 8639 3238
rect 10374 6010 10430 6012
rect 10454 6010 10510 6012
rect 10534 6010 10590 6012
rect 10614 6010 10670 6012
rect 10374 5958 10420 6010
rect 10420 5958 10430 6010
rect 10454 5958 10484 6010
rect 10484 5958 10496 6010
rect 10496 5958 10510 6010
rect 10534 5958 10548 6010
rect 10548 5958 10560 6010
rect 10560 5958 10590 6010
rect 10614 5958 10624 6010
rect 10624 5958 10670 6010
rect 10374 5956 10430 5958
rect 10454 5956 10510 5958
rect 10534 5956 10590 5958
rect 10614 5956 10670 5958
rect 10374 4922 10430 4924
rect 10454 4922 10510 4924
rect 10534 4922 10590 4924
rect 10614 4922 10670 4924
rect 10374 4870 10420 4922
rect 10420 4870 10430 4922
rect 10454 4870 10484 4922
rect 10484 4870 10496 4922
rect 10496 4870 10510 4922
rect 10534 4870 10548 4922
rect 10548 4870 10560 4922
rect 10560 4870 10590 4922
rect 10614 4870 10624 4922
rect 10624 4870 10670 4922
rect 10374 4868 10430 4870
rect 10454 4868 10510 4870
rect 10534 4868 10590 4870
rect 10614 4868 10670 4870
rect 10374 3834 10430 3836
rect 10454 3834 10510 3836
rect 10534 3834 10590 3836
rect 10614 3834 10670 3836
rect 10374 3782 10420 3834
rect 10420 3782 10430 3834
rect 10454 3782 10484 3834
rect 10484 3782 10496 3834
rect 10496 3782 10510 3834
rect 10534 3782 10548 3834
rect 10548 3782 10560 3834
rect 10560 3782 10590 3834
rect 10614 3782 10624 3834
rect 10624 3782 10670 3834
rect 10374 3780 10430 3782
rect 10454 3780 10510 3782
rect 10534 3780 10590 3782
rect 10614 3780 10670 3782
rect 10374 2746 10430 2748
rect 10454 2746 10510 2748
rect 10534 2746 10590 2748
rect 10614 2746 10670 2748
rect 10374 2694 10420 2746
rect 10420 2694 10430 2746
rect 10454 2694 10484 2746
rect 10484 2694 10496 2746
rect 10496 2694 10510 2746
rect 10534 2694 10548 2746
rect 10548 2694 10560 2746
rect 10560 2694 10590 2746
rect 10614 2694 10624 2746
rect 10624 2694 10670 2746
rect 10374 2692 10430 2694
rect 10454 2692 10510 2694
rect 10534 2692 10590 2694
rect 10614 2692 10670 2694
rect 5652 2202 5708 2204
rect 5732 2202 5788 2204
rect 5812 2202 5868 2204
rect 5892 2202 5948 2204
rect 5652 2150 5698 2202
rect 5698 2150 5708 2202
rect 5732 2150 5762 2202
rect 5762 2150 5774 2202
rect 5774 2150 5788 2202
rect 5812 2150 5826 2202
rect 5826 2150 5838 2202
rect 5838 2150 5868 2202
rect 5892 2150 5902 2202
rect 5902 2150 5948 2202
rect 5652 2148 5708 2150
rect 5732 2148 5788 2150
rect 5812 2148 5868 2150
rect 5892 2148 5948 2150
rect 8343 2202 8399 2204
rect 8423 2202 8479 2204
rect 8503 2202 8559 2204
rect 8583 2202 8639 2204
rect 8343 2150 8389 2202
rect 8389 2150 8399 2202
rect 8423 2150 8453 2202
rect 8453 2150 8465 2202
rect 8465 2150 8479 2202
rect 8503 2150 8517 2202
rect 8517 2150 8529 2202
rect 8529 2150 8559 2202
rect 8583 2150 8593 2202
rect 8593 2150 8639 2202
rect 8343 2148 8399 2150
rect 8423 2148 8479 2150
rect 8503 2148 8559 2150
rect 8583 2148 8639 2150
rect 11034 7642 11090 7644
rect 11114 7642 11170 7644
rect 11194 7642 11250 7644
rect 11274 7642 11330 7644
rect 11034 7590 11080 7642
rect 11080 7590 11090 7642
rect 11114 7590 11144 7642
rect 11144 7590 11156 7642
rect 11156 7590 11170 7642
rect 11194 7590 11208 7642
rect 11208 7590 11220 7642
rect 11220 7590 11250 7642
rect 11274 7590 11284 7642
rect 11284 7590 11330 7642
rect 11034 7588 11090 7590
rect 11114 7588 11170 7590
rect 11194 7588 11250 7590
rect 11274 7588 11330 7590
rect 11034 6554 11090 6556
rect 11114 6554 11170 6556
rect 11194 6554 11250 6556
rect 11274 6554 11330 6556
rect 11034 6502 11080 6554
rect 11080 6502 11090 6554
rect 11114 6502 11144 6554
rect 11144 6502 11156 6554
rect 11156 6502 11170 6554
rect 11194 6502 11208 6554
rect 11208 6502 11220 6554
rect 11220 6502 11250 6554
rect 11274 6502 11284 6554
rect 11284 6502 11330 6554
rect 11034 6500 11090 6502
rect 11114 6500 11170 6502
rect 11194 6500 11250 6502
rect 11274 6500 11330 6502
rect 11794 6160 11850 6216
rect 11034 5466 11090 5468
rect 11114 5466 11170 5468
rect 11194 5466 11250 5468
rect 11274 5466 11330 5468
rect 11034 5414 11080 5466
rect 11080 5414 11090 5466
rect 11114 5414 11144 5466
rect 11144 5414 11156 5466
rect 11156 5414 11170 5466
rect 11194 5414 11208 5466
rect 11208 5414 11220 5466
rect 11220 5414 11250 5466
rect 11274 5414 11284 5466
rect 11284 5414 11330 5466
rect 11034 5412 11090 5414
rect 11114 5412 11170 5414
rect 11194 5412 11250 5414
rect 11274 5412 11330 5414
rect 11034 4378 11090 4380
rect 11114 4378 11170 4380
rect 11194 4378 11250 4380
rect 11274 4378 11330 4380
rect 11034 4326 11080 4378
rect 11080 4326 11090 4378
rect 11114 4326 11144 4378
rect 11144 4326 11156 4378
rect 11156 4326 11170 4378
rect 11194 4326 11208 4378
rect 11208 4326 11220 4378
rect 11220 4326 11250 4378
rect 11274 4326 11284 4378
rect 11284 4326 11330 4378
rect 11034 4324 11090 4326
rect 11114 4324 11170 4326
rect 11194 4324 11250 4326
rect 11274 4324 11330 4326
rect 11034 3290 11090 3292
rect 11114 3290 11170 3292
rect 11194 3290 11250 3292
rect 11274 3290 11330 3292
rect 11034 3238 11080 3290
rect 11080 3238 11090 3290
rect 11114 3238 11144 3290
rect 11144 3238 11156 3290
rect 11156 3238 11170 3290
rect 11194 3238 11208 3290
rect 11208 3238 11220 3290
rect 11220 3238 11250 3290
rect 11274 3238 11284 3290
rect 11284 3238 11330 3290
rect 11034 3236 11090 3238
rect 11114 3236 11170 3238
rect 11194 3236 11250 3238
rect 11274 3236 11330 3238
rect 11034 2202 11090 2204
rect 11114 2202 11170 2204
rect 11194 2202 11250 2204
rect 11274 2202 11330 2204
rect 11034 2150 11080 2202
rect 11080 2150 11090 2202
rect 11114 2150 11144 2202
rect 11144 2150 11156 2202
rect 11156 2150 11170 2202
rect 11194 2150 11208 2202
rect 11208 2150 11220 2202
rect 11220 2150 11250 2202
rect 11274 2150 11284 2202
rect 11284 2150 11330 2202
rect 11034 2148 11090 2150
rect 11114 2148 11170 2150
rect 11194 2148 11250 2150
rect 11274 2148 11330 2150
rect 10874 720 10930 776
<< metal3 >>
rect 0 14378 800 14408
rect 0 14318 1042 14378
rect 0 14288 800 14318
rect 982 14106 1042 14318
rect 1393 14106 1459 14109
rect 982 14104 1459 14106
rect 982 14048 1398 14104
rect 1454 14048 1459 14104
rect 982 14046 1459 14048
rect 1393 14043 1459 14046
rect 2291 12544 2607 12545
rect 2291 12480 2297 12544
rect 2361 12480 2377 12544
rect 2441 12480 2457 12544
rect 2521 12480 2537 12544
rect 2601 12480 2607 12544
rect 2291 12479 2607 12480
rect 4982 12544 5298 12545
rect 4982 12480 4988 12544
rect 5052 12480 5068 12544
rect 5132 12480 5148 12544
rect 5212 12480 5228 12544
rect 5292 12480 5298 12544
rect 4982 12479 5298 12480
rect 7673 12544 7989 12545
rect 7673 12480 7679 12544
rect 7743 12480 7759 12544
rect 7823 12480 7839 12544
rect 7903 12480 7919 12544
rect 7983 12480 7989 12544
rect 7673 12479 7989 12480
rect 10364 12544 10680 12545
rect 10364 12480 10370 12544
rect 10434 12480 10450 12544
rect 10514 12480 10530 12544
rect 10594 12480 10610 12544
rect 10674 12480 10680 12544
rect 10364 12479 10680 12480
rect 11237 12338 11303 12341
rect 12202 12338 13002 12368
rect 11237 12336 13002 12338
rect 11237 12280 11242 12336
rect 11298 12280 13002 12336
rect 11237 12278 13002 12280
rect 11237 12275 11303 12278
rect 12202 12248 13002 12278
rect 2951 12000 3267 12001
rect 2951 11936 2957 12000
rect 3021 11936 3037 12000
rect 3101 11936 3117 12000
rect 3181 11936 3197 12000
rect 3261 11936 3267 12000
rect 2951 11935 3267 11936
rect 5642 12000 5958 12001
rect 5642 11936 5648 12000
rect 5712 11936 5728 12000
rect 5792 11936 5808 12000
rect 5872 11936 5888 12000
rect 5952 11936 5958 12000
rect 5642 11935 5958 11936
rect 8333 12000 8649 12001
rect 8333 11936 8339 12000
rect 8403 11936 8419 12000
rect 8483 11936 8499 12000
rect 8563 11936 8579 12000
rect 8643 11936 8649 12000
rect 8333 11935 8649 11936
rect 11024 12000 11340 12001
rect 11024 11936 11030 12000
rect 11094 11936 11110 12000
rect 11174 11936 11190 12000
rect 11254 11936 11270 12000
rect 11334 11936 11340 12000
rect 11024 11935 11340 11936
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 2291 11456 2607 11457
rect 2291 11392 2297 11456
rect 2361 11392 2377 11456
rect 2441 11392 2457 11456
rect 2521 11392 2537 11456
rect 2601 11392 2607 11456
rect 2291 11391 2607 11392
rect 4982 11456 5298 11457
rect 4982 11392 4988 11456
rect 5052 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5298 11456
rect 4982 11391 5298 11392
rect 7673 11456 7989 11457
rect 7673 11392 7679 11456
rect 7743 11392 7759 11456
rect 7823 11392 7839 11456
rect 7903 11392 7919 11456
rect 7983 11392 7989 11456
rect 7673 11391 7989 11392
rect 10364 11456 10680 11457
rect 10364 11392 10370 11456
rect 10434 11392 10450 11456
rect 10514 11392 10530 11456
rect 10594 11392 10610 11456
rect 10674 11392 10680 11456
rect 10364 11391 10680 11392
rect 2951 10912 3267 10913
rect 2951 10848 2957 10912
rect 3021 10848 3037 10912
rect 3101 10848 3117 10912
rect 3181 10848 3197 10912
rect 3261 10848 3267 10912
rect 2951 10847 3267 10848
rect 5642 10912 5958 10913
rect 5642 10848 5648 10912
rect 5712 10848 5728 10912
rect 5792 10848 5808 10912
rect 5872 10848 5888 10912
rect 5952 10848 5958 10912
rect 5642 10847 5958 10848
rect 8333 10912 8649 10913
rect 8333 10848 8339 10912
rect 8403 10848 8419 10912
rect 8483 10848 8499 10912
rect 8563 10848 8579 10912
rect 8643 10848 8649 10912
rect 8333 10847 8649 10848
rect 11024 10912 11340 10913
rect 11024 10848 11030 10912
rect 11094 10848 11110 10912
rect 11174 10848 11190 10912
rect 11254 10848 11270 10912
rect 11334 10848 11340 10912
rect 11024 10847 11340 10848
rect 2497 10706 2563 10709
rect 5441 10706 5507 10709
rect 2497 10704 5507 10706
rect 2497 10648 2502 10704
rect 2558 10648 5446 10704
rect 5502 10648 5507 10704
rect 2497 10646 5507 10648
rect 2497 10643 2563 10646
rect 5441 10643 5507 10646
rect 2291 10368 2607 10369
rect 2291 10304 2297 10368
rect 2361 10304 2377 10368
rect 2441 10304 2457 10368
rect 2521 10304 2537 10368
rect 2601 10304 2607 10368
rect 2291 10303 2607 10304
rect 4982 10368 5298 10369
rect 4982 10304 4988 10368
rect 5052 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5298 10368
rect 4982 10303 5298 10304
rect 7673 10368 7989 10369
rect 7673 10304 7679 10368
rect 7743 10304 7759 10368
rect 7823 10304 7839 10368
rect 7903 10304 7919 10368
rect 7983 10304 7989 10368
rect 7673 10303 7989 10304
rect 10364 10368 10680 10369
rect 10364 10304 10370 10368
rect 10434 10304 10450 10368
rect 10514 10304 10530 10368
rect 10594 10304 10610 10368
rect 10674 10304 10680 10368
rect 10364 10303 10680 10304
rect 2951 9824 3267 9825
rect 2951 9760 2957 9824
rect 3021 9760 3037 9824
rect 3101 9760 3117 9824
rect 3181 9760 3197 9824
rect 3261 9760 3267 9824
rect 2951 9759 3267 9760
rect 5642 9824 5958 9825
rect 5642 9760 5648 9824
rect 5712 9760 5728 9824
rect 5792 9760 5808 9824
rect 5872 9760 5888 9824
rect 5952 9760 5958 9824
rect 5642 9759 5958 9760
rect 8333 9824 8649 9825
rect 8333 9760 8339 9824
rect 8403 9760 8419 9824
rect 8483 9760 8499 9824
rect 8563 9760 8579 9824
rect 8643 9760 8649 9824
rect 8333 9759 8649 9760
rect 11024 9824 11340 9825
rect 11024 9760 11030 9824
rect 11094 9760 11110 9824
rect 11174 9760 11190 9824
rect 11254 9760 11270 9824
rect 11334 9760 11340 9824
rect 11024 9759 11340 9760
rect 12065 9618 12131 9621
rect 12202 9618 13002 9648
rect 12065 9616 13002 9618
rect 12065 9560 12070 9616
rect 12126 9560 13002 9616
rect 12065 9558 13002 9560
rect 12065 9555 12131 9558
rect 12202 9528 13002 9558
rect 2291 9280 2607 9281
rect 2291 9216 2297 9280
rect 2361 9216 2377 9280
rect 2441 9216 2457 9280
rect 2521 9216 2537 9280
rect 2601 9216 2607 9280
rect 2291 9215 2607 9216
rect 4982 9280 5298 9281
rect 4982 9216 4988 9280
rect 5052 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5298 9280
rect 4982 9215 5298 9216
rect 7673 9280 7989 9281
rect 7673 9216 7679 9280
rect 7743 9216 7759 9280
rect 7823 9216 7839 9280
rect 7903 9216 7919 9280
rect 7983 9216 7989 9280
rect 7673 9215 7989 9216
rect 10364 9280 10680 9281
rect 10364 9216 10370 9280
rect 10434 9216 10450 9280
rect 10514 9216 10530 9280
rect 10594 9216 10610 9280
rect 10674 9216 10680 9280
rect 10364 9215 10680 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 2951 8736 3267 8737
rect 2951 8672 2957 8736
rect 3021 8672 3037 8736
rect 3101 8672 3117 8736
rect 3181 8672 3197 8736
rect 3261 8672 3267 8736
rect 2951 8671 3267 8672
rect 5642 8736 5958 8737
rect 5642 8672 5648 8736
rect 5712 8672 5728 8736
rect 5792 8672 5808 8736
rect 5872 8672 5888 8736
rect 5952 8672 5958 8736
rect 5642 8671 5958 8672
rect 8333 8736 8649 8737
rect 8333 8672 8339 8736
rect 8403 8672 8419 8736
rect 8483 8672 8499 8736
rect 8563 8672 8579 8736
rect 8643 8672 8649 8736
rect 8333 8671 8649 8672
rect 11024 8736 11340 8737
rect 11024 8672 11030 8736
rect 11094 8672 11110 8736
rect 11174 8672 11190 8736
rect 11254 8672 11270 8736
rect 11334 8672 11340 8736
rect 11024 8671 11340 8672
rect 2291 8192 2607 8193
rect 2291 8128 2297 8192
rect 2361 8128 2377 8192
rect 2441 8128 2457 8192
rect 2521 8128 2537 8192
rect 2601 8128 2607 8192
rect 2291 8127 2607 8128
rect 4982 8192 5298 8193
rect 4982 8128 4988 8192
rect 5052 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5298 8192
rect 4982 8127 5298 8128
rect 7673 8192 7989 8193
rect 7673 8128 7679 8192
rect 7743 8128 7759 8192
rect 7823 8128 7839 8192
rect 7903 8128 7919 8192
rect 7983 8128 7989 8192
rect 7673 8127 7989 8128
rect 10364 8192 10680 8193
rect 10364 8128 10370 8192
rect 10434 8128 10450 8192
rect 10514 8128 10530 8192
rect 10594 8128 10610 8192
rect 10674 8128 10680 8192
rect 10364 8127 10680 8128
rect 2951 7648 3267 7649
rect 2951 7584 2957 7648
rect 3021 7584 3037 7648
rect 3101 7584 3117 7648
rect 3181 7584 3197 7648
rect 3261 7584 3267 7648
rect 2951 7583 3267 7584
rect 5642 7648 5958 7649
rect 5642 7584 5648 7648
rect 5712 7584 5728 7648
rect 5792 7584 5808 7648
rect 5872 7584 5888 7648
rect 5952 7584 5958 7648
rect 5642 7583 5958 7584
rect 8333 7648 8649 7649
rect 8333 7584 8339 7648
rect 8403 7584 8419 7648
rect 8483 7584 8499 7648
rect 8563 7584 8579 7648
rect 8643 7584 8649 7648
rect 8333 7583 8649 7584
rect 11024 7648 11340 7649
rect 11024 7584 11030 7648
rect 11094 7584 11110 7648
rect 11174 7584 11190 7648
rect 11254 7584 11270 7648
rect 11334 7584 11340 7648
rect 11024 7583 11340 7584
rect 2291 7104 2607 7105
rect 2291 7040 2297 7104
rect 2361 7040 2377 7104
rect 2441 7040 2457 7104
rect 2521 7040 2537 7104
rect 2601 7040 2607 7104
rect 2291 7039 2607 7040
rect 4982 7104 5298 7105
rect 4982 7040 4988 7104
rect 5052 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5298 7104
rect 4982 7039 5298 7040
rect 7673 7104 7989 7105
rect 7673 7040 7679 7104
rect 7743 7040 7759 7104
rect 7823 7040 7839 7104
rect 7903 7040 7919 7104
rect 7983 7040 7989 7104
rect 7673 7039 7989 7040
rect 10364 7104 10680 7105
rect 10364 7040 10370 7104
rect 10434 7040 10450 7104
rect 10514 7040 10530 7104
rect 10594 7040 10610 7104
rect 10674 7040 10680 7104
rect 10364 7039 10680 7040
rect 6913 7036 6979 7037
rect 6862 6972 6868 7036
rect 6932 7034 6979 7036
rect 8201 7034 8267 7037
rect 9622 7034 9628 7036
rect 6932 7032 7024 7034
rect 6974 6976 7024 7032
rect 6932 6974 7024 6976
rect 8201 7032 9628 7034
rect 8201 6976 8206 7032
rect 8262 6976 9628 7032
rect 8201 6974 9628 6976
rect 6932 6972 6979 6974
rect 6913 6971 6979 6972
rect 8201 6971 8267 6974
rect 9622 6972 9628 6974
rect 9692 6972 9698 7036
rect 6269 6762 6335 6765
rect 7557 6762 7623 6765
rect 6269 6760 7623 6762
rect 6269 6704 6274 6760
rect 6330 6704 7562 6760
rect 7618 6704 7623 6760
rect 6269 6702 7623 6704
rect 6269 6699 6335 6702
rect 7557 6699 7623 6702
rect 2951 6560 3267 6561
rect 2951 6496 2957 6560
rect 3021 6496 3037 6560
rect 3101 6496 3117 6560
rect 3181 6496 3197 6560
rect 3261 6496 3267 6560
rect 2951 6495 3267 6496
rect 5642 6560 5958 6561
rect 5642 6496 5648 6560
rect 5712 6496 5728 6560
rect 5792 6496 5808 6560
rect 5872 6496 5888 6560
rect 5952 6496 5958 6560
rect 5642 6495 5958 6496
rect 8333 6560 8649 6561
rect 8333 6496 8339 6560
rect 8403 6496 8419 6560
rect 8483 6496 8499 6560
rect 8563 6496 8579 6560
rect 8643 6496 8649 6560
rect 8333 6495 8649 6496
rect 11024 6560 11340 6561
rect 11024 6496 11030 6560
rect 11094 6496 11110 6560
rect 11174 6496 11190 6560
rect 11254 6496 11270 6560
rect 11334 6496 11340 6560
rect 11024 6495 11340 6496
rect 6913 6354 6979 6357
rect 9029 6354 9095 6357
rect 6913 6352 9095 6354
rect 6913 6296 6918 6352
rect 6974 6296 9034 6352
rect 9090 6296 9095 6352
rect 6913 6294 9095 6296
rect 6913 6291 6979 6294
rect 9029 6291 9095 6294
rect 11789 6218 11855 6221
rect 12202 6218 13002 6248
rect 11789 6216 13002 6218
rect 11789 6160 11794 6216
rect 11850 6160 13002 6216
rect 11789 6158 13002 6160
rect 11789 6155 11855 6158
rect 12202 6128 13002 6158
rect 2291 6016 2607 6017
rect 2291 5952 2297 6016
rect 2361 5952 2377 6016
rect 2441 5952 2457 6016
rect 2521 5952 2537 6016
rect 2601 5952 2607 6016
rect 2291 5951 2607 5952
rect 4982 6016 5298 6017
rect 4982 5952 4988 6016
rect 5052 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5298 6016
rect 4982 5951 5298 5952
rect 7673 6016 7989 6017
rect 7673 5952 7679 6016
rect 7743 5952 7759 6016
rect 7823 5952 7839 6016
rect 7903 5952 7919 6016
rect 7983 5952 7989 6016
rect 7673 5951 7989 5952
rect 10364 6016 10680 6017
rect 10364 5952 10370 6016
rect 10434 5952 10450 6016
rect 10514 5952 10530 6016
rect 10594 5952 10610 6016
rect 10674 5952 10680 6016
rect 10364 5951 10680 5952
rect 0 5538 800 5568
rect 933 5538 999 5541
rect 0 5536 999 5538
rect 0 5480 938 5536
rect 994 5480 999 5536
rect 0 5478 999 5480
rect 0 5448 800 5478
rect 933 5475 999 5478
rect 2951 5472 3267 5473
rect 2951 5408 2957 5472
rect 3021 5408 3037 5472
rect 3101 5408 3117 5472
rect 3181 5408 3197 5472
rect 3261 5408 3267 5472
rect 2951 5407 3267 5408
rect 5642 5472 5958 5473
rect 5642 5408 5648 5472
rect 5712 5408 5728 5472
rect 5792 5408 5808 5472
rect 5872 5408 5888 5472
rect 5952 5408 5958 5472
rect 5642 5407 5958 5408
rect 8333 5472 8649 5473
rect 8333 5408 8339 5472
rect 8403 5408 8419 5472
rect 8483 5408 8499 5472
rect 8563 5408 8579 5472
rect 8643 5408 8649 5472
rect 8333 5407 8649 5408
rect 11024 5472 11340 5473
rect 11024 5408 11030 5472
rect 11094 5408 11110 5472
rect 11174 5408 11190 5472
rect 11254 5408 11270 5472
rect 11334 5408 11340 5472
rect 11024 5407 11340 5408
rect 2291 4928 2607 4929
rect 2291 4864 2297 4928
rect 2361 4864 2377 4928
rect 2441 4864 2457 4928
rect 2521 4864 2537 4928
rect 2601 4864 2607 4928
rect 2291 4863 2607 4864
rect 4982 4928 5298 4929
rect 4982 4864 4988 4928
rect 5052 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5298 4928
rect 4982 4863 5298 4864
rect 7673 4928 7989 4929
rect 7673 4864 7679 4928
rect 7743 4864 7759 4928
rect 7823 4864 7839 4928
rect 7903 4864 7919 4928
rect 7983 4864 7989 4928
rect 7673 4863 7989 4864
rect 10364 4928 10680 4929
rect 10364 4864 10370 4928
rect 10434 4864 10450 4928
rect 10514 4864 10530 4928
rect 10594 4864 10610 4928
rect 10674 4864 10680 4928
rect 10364 4863 10680 4864
rect 2951 4384 3267 4385
rect 2951 4320 2957 4384
rect 3021 4320 3037 4384
rect 3101 4320 3117 4384
rect 3181 4320 3197 4384
rect 3261 4320 3267 4384
rect 2951 4319 3267 4320
rect 5642 4384 5958 4385
rect 5642 4320 5648 4384
rect 5712 4320 5728 4384
rect 5792 4320 5808 4384
rect 5872 4320 5888 4384
rect 5952 4320 5958 4384
rect 5642 4319 5958 4320
rect 8333 4384 8649 4385
rect 8333 4320 8339 4384
rect 8403 4320 8419 4384
rect 8483 4320 8499 4384
rect 8563 4320 8579 4384
rect 8643 4320 8649 4384
rect 8333 4319 8649 4320
rect 11024 4384 11340 4385
rect 11024 4320 11030 4384
rect 11094 4320 11110 4384
rect 11174 4320 11190 4384
rect 11254 4320 11270 4384
rect 11334 4320 11340 4384
rect 11024 4319 11340 4320
rect 6177 4042 6243 4045
rect 6862 4042 6868 4044
rect 6177 4040 6868 4042
rect 6177 3984 6182 4040
rect 6238 3984 6868 4040
rect 6177 3982 6868 3984
rect 6177 3979 6243 3982
rect 6862 3980 6868 3982
rect 6932 3980 6938 4044
rect 2291 3840 2607 3841
rect 2291 3776 2297 3840
rect 2361 3776 2377 3840
rect 2441 3776 2457 3840
rect 2521 3776 2537 3840
rect 2601 3776 2607 3840
rect 2291 3775 2607 3776
rect 4982 3840 5298 3841
rect 4982 3776 4988 3840
rect 5052 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5298 3840
rect 4982 3775 5298 3776
rect 7673 3840 7989 3841
rect 7673 3776 7679 3840
rect 7743 3776 7759 3840
rect 7823 3776 7839 3840
rect 7903 3776 7919 3840
rect 7983 3776 7989 3840
rect 7673 3775 7989 3776
rect 10364 3840 10680 3841
rect 10364 3776 10370 3840
rect 10434 3776 10450 3840
rect 10514 3776 10530 3840
rect 10594 3776 10610 3840
rect 10674 3776 10680 3840
rect 10364 3775 10680 3776
rect 9622 3436 9628 3500
rect 9692 3498 9698 3500
rect 12202 3498 13002 3528
rect 9692 3438 13002 3498
rect 9692 3436 9698 3438
rect 12202 3408 13002 3438
rect 2951 3296 3267 3297
rect 2951 3232 2957 3296
rect 3021 3232 3037 3296
rect 3101 3232 3117 3296
rect 3181 3232 3197 3296
rect 3261 3232 3267 3296
rect 2951 3231 3267 3232
rect 5642 3296 5958 3297
rect 5642 3232 5648 3296
rect 5712 3232 5728 3296
rect 5792 3232 5808 3296
rect 5872 3232 5888 3296
rect 5952 3232 5958 3296
rect 5642 3231 5958 3232
rect 8333 3296 8649 3297
rect 8333 3232 8339 3296
rect 8403 3232 8419 3296
rect 8483 3232 8499 3296
rect 8563 3232 8579 3296
rect 8643 3232 8649 3296
rect 8333 3231 8649 3232
rect 11024 3296 11340 3297
rect 11024 3232 11030 3296
rect 11094 3232 11110 3296
rect 11174 3232 11190 3296
rect 11254 3232 11270 3296
rect 11334 3232 11340 3296
rect 11024 3231 11340 3232
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 2291 2752 2607 2753
rect 2291 2688 2297 2752
rect 2361 2688 2377 2752
rect 2441 2688 2457 2752
rect 2521 2688 2537 2752
rect 2601 2688 2607 2752
rect 2291 2687 2607 2688
rect 4982 2752 5298 2753
rect 4982 2688 4988 2752
rect 5052 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5298 2752
rect 4982 2687 5298 2688
rect 7673 2752 7989 2753
rect 7673 2688 7679 2752
rect 7743 2688 7759 2752
rect 7823 2688 7839 2752
rect 7903 2688 7919 2752
rect 7983 2688 7989 2752
rect 7673 2687 7989 2688
rect 10364 2752 10680 2753
rect 10364 2688 10370 2752
rect 10434 2688 10450 2752
rect 10514 2688 10530 2752
rect 10594 2688 10610 2752
rect 10674 2688 10680 2752
rect 10364 2687 10680 2688
rect 2951 2208 3267 2209
rect 2951 2144 2957 2208
rect 3021 2144 3037 2208
rect 3101 2144 3117 2208
rect 3181 2144 3197 2208
rect 3261 2144 3267 2208
rect 2951 2143 3267 2144
rect 5642 2208 5958 2209
rect 5642 2144 5648 2208
rect 5712 2144 5728 2208
rect 5792 2144 5808 2208
rect 5872 2144 5888 2208
rect 5952 2144 5958 2208
rect 5642 2143 5958 2144
rect 8333 2208 8649 2209
rect 8333 2144 8339 2208
rect 8403 2144 8419 2208
rect 8483 2144 8499 2208
rect 8563 2144 8579 2208
rect 8643 2144 8649 2208
rect 8333 2143 8649 2144
rect 11024 2208 11340 2209
rect 11024 2144 11030 2208
rect 11094 2144 11110 2208
rect 11174 2144 11190 2208
rect 11254 2144 11270 2208
rect 11334 2144 11340 2208
rect 11024 2143 11340 2144
rect 10869 778 10935 781
rect 12202 778 13002 808
rect 10869 776 13002 778
rect 10869 720 10874 776
rect 10930 720 13002 776
rect 10869 718 13002 720
rect 10869 715 10935 718
rect 12202 688 13002 718
<< via3 >>
rect 2297 12540 2361 12544
rect 2297 12484 2301 12540
rect 2301 12484 2357 12540
rect 2357 12484 2361 12540
rect 2297 12480 2361 12484
rect 2377 12540 2441 12544
rect 2377 12484 2381 12540
rect 2381 12484 2437 12540
rect 2437 12484 2441 12540
rect 2377 12480 2441 12484
rect 2457 12540 2521 12544
rect 2457 12484 2461 12540
rect 2461 12484 2517 12540
rect 2517 12484 2521 12540
rect 2457 12480 2521 12484
rect 2537 12540 2601 12544
rect 2537 12484 2541 12540
rect 2541 12484 2597 12540
rect 2597 12484 2601 12540
rect 2537 12480 2601 12484
rect 4988 12540 5052 12544
rect 4988 12484 4992 12540
rect 4992 12484 5048 12540
rect 5048 12484 5052 12540
rect 4988 12480 5052 12484
rect 5068 12540 5132 12544
rect 5068 12484 5072 12540
rect 5072 12484 5128 12540
rect 5128 12484 5132 12540
rect 5068 12480 5132 12484
rect 5148 12540 5212 12544
rect 5148 12484 5152 12540
rect 5152 12484 5208 12540
rect 5208 12484 5212 12540
rect 5148 12480 5212 12484
rect 5228 12540 5292 12544
rect 5228 12484 5232 12540
rect 5232 12484 5288 12540
rect 5288 12484 5292 12540
rect 5228 12480 5292 12484
rect 7679 12540 7743 12544
rect 7679 12484 7683 12540
rect 7683 12484 7739 12540
rect 7739 12484 7743 12540
rect 7679 12480 7743 12484
rect 7759 12540 7823 12544
rect 7759 12484 7763 12540
rect 7763 12484 7819 12540
rect 7819 12484 7823 12540
rect 7759 12480 7823 12484
rect 7839 12540 7903 12544
rect 7839 12484 7843 12540
rect 7843 12484 7899 12540
rect 7899 12484 7903 12540
rect 7839 12480 7903 12484
rect 7919 12540 7983 12544
rect 7919 12484 7923 12540
rect 7923 12484 7979 12540
rect 7979 12484 7983 12540
rect 7919 12480 7983 12484
rect 10370 12540 10434 12544
rect 10370 12484 10374 12540
rect 10374 12484 10430 12540
rect 10430 12484 10434 12540
rect 10370 12480 10434 12484
rect 10450 12540 10514 12544
rect 10450 12484 10454 12540
rect 10454 12484 10510 12540
rect 10510 12484 10514 12540
rect 10450 12480 10514 12484
rect 10530 12540 10594 12544
rect 10530 12484 10534 12540
rect 10534 12484 10590 12540
rect 10590 12484 10594 12540
rect 10530 12480 10594 12484
rect 10610 12540 10674 12544
rect 10610 12484 10614 12540
rect 10614 12484 10670 12540
rect 10670 12484 10674 12540
rect 10610 12480 10674 12484
rect 2957 11996 3021 12000
rect 2957 11940 2961 11996
rect 2961 11940 3017 11996
rect 3017 11940 3021 11996
rect 2957 11936 3021 11940
rect 3037 11996 3101 12000
rect 3037 11940 3041 11996
rect 3041 11940 3097 11996
rect 3097 11940 3101 11996
rect 3037 11936 3101 11940
rect 3117 11996 3181 12000
rect 3117 11940 3121 11996
rect 3121 11940 3177 11996
rect 3177 11940 3181 11996
rect 3117 11936 3181 11940
rect 3197 11996 3261 12000
rect 3197 11940 3201 11996
rect 3201 11940 3257 11996
rect 3257 11940 3261 11996
rect 3197 11936 3261 11940
rect 5648 11996 5712 12000
rect 5648 11940 5652 11996
rect 5652 11940 5708 11996
rect 5708 11940 5712 11996
rect 5648 11936 5712 11940
rect 5728 11996 5792 12000
rect 5728 11940 5732 11996
rect 5732 11940 5788 11996
rect 5788 11940 5792 11996
rect 5728 11936 5792 11940
rect 5808 11996 5872 12000
rect 5808 11940 5812 11996
rect 5812 11940 5868 11996
rect 5868 11940 5872 11996
rect 5808 11936 5872 11940
rect 5888 11996 5952 12000
rect 5888 11940 5892 11996
rect 5892 11940 5948 11996
rect 5948 11940 5952 11996
rect 5888 11936 5952 11940
rect 8339 11996 8403 12000
rect 8339 11940 8343 11996
rect 8343 11940 8399 11996
rect 8399 11940 8403 11996
rect 8339 11936 8403 11940
rect 8419 11996 8483 12000
rect 8419 11940 8423 11996
rect 8423 11940 8479 11996
rect 8479 11940 8483 11996
rect 8419 11936 8483 11940
rect 8499 11996 8563 12000
rect 8499 11940 8503 11996
rect 8503 11940 8559 11996
rect 8559 11940 8563 11996
rect 8499 11936 8563 11940
rect 8579 11996 8643 12000
rect 8579 11940 8583 11996
rect 8583 11940 8639 11996
rect 8639 11940 8643 11996
rect 8579 11936 8643 11940
rect 11030 11996 11094 12000
rect 11030 11940 11034 11996
rect 11034 11940 11090 11996
rect 11090 11940 11094 11996
rect 11030 11936 11094 11940
rect 11110 11996 11174 12000
rect 11110 11940 11114 11996
rect 11114 11940 11170 11996
rect 11170 11940 11174 11996
rect 11110 11936 11174 11940
rect 11190 11996 11254 12000
rect 11190 11940 11194 11996
rect 11194 11940 11250 11996
rect 11250 11940 11254 11996
rect 11190 11936 11254 11940
rect 11270 11996 11334 12000
rect 11270 11940 11274 11996
rect 11274 11940 11330 11996
rect 11330 11940 11334 11996
rect 11270 11936 11334 11940
rect 2297 11452 2361 11456
rect 2297 11396 2301 11452
rect 2301 11396 2357 11452
rect 2357 11396 2361 11452
rect 2297 11392 2361 11396
rect 2377 11452 2441 11456
rect 2377 11396 2381 11452
rect 2381 11396 2437 11452
rect 2437 11396 2441 11452
rect 2377 11392 2441 11396
rect 2457 11452 2521 11456
rect 2457 11396 2461 11452
rect 2461 11396 2517 11452
rect 2517 11396 2521 11452
rect 2457 11392 2521 11396
rect 2537 11452 2601 11456
rect 2537 11396 2541 11452
rect 2541 11396 2597 11452
rect 2597 11396 2601 11452
rect 2537 11392 2601 11396
rect 4988 11452 5052 11456
rect 4988 11396 4992 11452
rect 4992 11396 5048 11452
rect 5048 11396 5052 11452
rect 4988 11392 5052 11396
rect 5068 11452 5132 11456
rect 5068 11396 5072 11452
rect 5072 11396 5128 11452
rect 5128 11396 5132 11452
rect 5068 11392 5132 11396
rect 5148 11452 5212 11456
rect 5148 11396 5152 11452
rect 5152 11396 5208 11452
rect 5208 11396 5212 11452
rect 5148 11392 5212 11396
rect 5228 11452 5292 11456
rect 5228 11396 5232 11452
rect 5232 11396 5288 11452
rect 5288 11396 5292 11452
rect 5228 11392 5292 11396
rect 7679 11452 7743 11456
rect 7679 11396 7683 11452
rect 7683 11396 7739 11452
rect 7739 11396 7743 11452
rect 7679 11392 7743 11396
rect 7759 11452 7823 11456
rect 7759 11396 7763 11452
rect 7763 11396 7819 11452
rect 7819 11396 7823 11452
rect 7759 11392 7823 11396
rect 7839 11452 7903 11456
rect 7839 11396 7843 11452
rect 7843 11396 7899 11452
rect 7899 11396 7903 11452
rect 7839 11392 7903 11396
rect 7919 11452 7983 11456
rect 7919 11396 7923 11452
rect 7923 11396 7979 11452
rect 7979 11396 7983 11452
rect 7919 11392 7983 11396
rect 10370 11452 10434 11456
rect 10370 11396 10374 11452
rect 10374 11396 10430 11452
rect 10430 11396 10434 11452
rect 10370 11392 10434 11396
rect 10450 11452 10514 11456
rect 10450 11396 10454 11452
rect 10454 11396 10510 11452
rect 10510 11396 10514 11452
rect 10450 11392 10514 11396
rect 10530 11452 10594 11456
rect 10530 11396 10534 11452
rect 10534 11396 10590 11452
rect 10590 11396 10594 11452
rect 10530 11392 10594 11396
rect 10610 11452 10674 11456
rect 10610 11396 10614 11452
rect 10614 11396 10670 11452
rect 10670 11396 10674 11452
rect 10610 11392 10674 11396
rect 2957 10908 3021 10912
rect 2957 10852 2961 10908
rect 2961 10852 3017 10908
rect 3017 10852 3021 10908
rect 2957 10848 3021 10852
rect 3037 10908 3101 10912
rect 3037 10852 3041 10908
rect 3041 10852 3097 10908
rect 3097 10852 3101 10908
rect 3037 10848 3101 10852
rect 3117 10908 3181 10912
rect 3117 10852 3121 10908
rect 3121 10852 3177 10908
rect 3177 10852 3181 10908
rect 3117 10848 3181 10852
rect 3197 10908 3261 10912
rect 3197 10852 3201 10908
rect 3201 10852 3257 10908
rect 3257 10852 3261 10908
rect 3197 10848 3261 10852
rect 5648 10908 5712 10912
rect 5648 10852 5652 10908
rect 5652 10852 5708 10908
rect 5708 10852 5712 10908
rect 5648 10848 5712 10852
rect 5728 10908 5792 10912
rect 5728 10852 5732 10908
rect 5732 10852 5788 10908
rect 5788 10852 5792 10908
rect 5728 10848 5792 10852
rect 5808 10908 5872 10912
rect 5808 10852 5812 10908
rect 5812 10852 5868 10908
rect 5868 10852 5872 10908
rect 5808 10848 5872 10852
rect 5888 10908 5952 10912
rect 5888 10852 5892 10908
rect 5892 10852 5948 10908
rect 5948 10852 5952 10908
rect 5888 10848 5952 10852
rect 8339 10908 8403 10912
rect 8339 10852 8343 10908
rect 8343 10852 8399 10908
rect 8399 10852 8403 10908
rect 8339 10848 8403 10852
rect 8419 10908 8483 10912
rect 8419 10852 8423 10908
rect 8423 10852 8479 10908
rect 8479 10852 8483 10908
rect 8419 10848 8483 10852
rect 8499 10908 8563 10912
rect 8499 10852 8503 10908
rect 8503 10852 8559 10908
rect 8559 10852 8563 10908
rect 8499 10848 8563 10852
rect 8579 10908 8643 10912
rect 8579 10852 8583 10908
rect 8583 10852 8639 10908
rect 8639 10852 8643 10908
rect 8579 10848 8643 10852
rect 11030 10908 11094 10912
rect 11030 10852 11034 10908
rect 11034 10852 11090 10908
rect 11090 10852 11094 10908
rect 11030 10848 11094 10852
rect 11110 10908 11174 10912
rect 11110 10852 11114 10908
rect 11114 10852 11170 10908
rect 11170 10852 11174 10908
rect 11110 10848 11174 10852
rect 11190 10908 11254 10912
rect 11190 10852 11194 10908
rect 11194 10852 11250 10908
rect 11250 10852 11254 10908
rect 11190 10848 11254 10852
rect 11270 10908 11334 10912
rect 11270 10852 11274 10908
rect 11274 10852 11330 10908
rect 11330 10852 11334 10908
rect 11270 10848 11334 10852
rect 2297 10364 2361 10368
rect 2297 10308 2301 10364
rect 2301 10308 2357 10364
rect 2357 10308 2361 10364
rect 2297 10304 2361 10308
rect 2377 10364 2441 10368
rect 2377 10308 2381 10364
rect 2381 10308 2437 10364
rect 2437 10308 2441 10364
rect 2377 10304 2441 10308
rect 2457 10364 2521 10368
rect 2457 10308 2461 10364
rect 2461 10308 2517 10364
rect 2517 10308 2521 10364
rect 2457 10304 2521 10308
rect 2537 10364 2601 10368
rect 2537 10308 2541 10364
rect 2541 10308 2597 10364
rect 2597 10308 2601 10364
rect 2537 10304 2601 10308
rect 4988 10364 5052 10368
rect 4988 10308 4992 10364
rect 4992 10308 5048 10364
rect 5048 10308 5052 10364
rect 4988 10304 5052 10308
rect 5068 10364 5132 10368
rect 5068 10308 5072 10364
rect 5072 10308 5128 10364
rect 5128 10308 5132 10364
rect 5068 10304 5132 10308
rect 5148 10364 5212 10368
rect 5148 10308 5152 10364
rect 5152 10308 5208 10364
rect 5208 10308 5212 10364
rect 5148 10304 5212 10308
rect 5228 10364 5292 10368
rect 5228 10308 5232 10364
rect 5232 10308 5288 10364
rect 5288 10308 5292 10364
rect 5228 10304 5292 10308
rect 7679 10364 7743 10368
rect 7679 10308 7683 10364
rect 7683 10308 7739 10364
rect 7739 10308 7743 10364
rect 7679 10304 7743 10308
rect 7759 10364 7823 10368
rect 7759 10308 7763 10364
rect 7763 10308 7819 10364
rect 7819 10308 7823 10364
rect 7759 10304 7823 10308
rect 7839 10364 7903 10368
rect 7839 10308 7843 10364
rect 7843 10308 7899 10364
rect 7899 10308 7903 10364
rect 7839 10304 7903 10308
rect 7919 10364 7983 10368
rect 7919 10308 7923 10364
rect 7923 10308 7979 10364
rect 7979 10308 7983 10364
rect 7919 10304 7983 10308
rect 10370 10364 10434 10368
rect 10370 10308 10374 10364
rect 10374 10308 10430 10364
rect 10430 10308 10434 10364
rect 10370 10304 10434 10308
rect 10450 10364 10514 10368
rect 10450 10308 10454 10364
rect 10454 10308 10510 10364
rect 10510 10308 10514 10364
rect 10450 10304 10514 10308
rect 10530 10364 10594 10368
rect 10530 10308 10534 10364
rect 10534 10308 10590 10364
rect 10590 10308 10594 10364
rect 10530 10304 10594 10308
rect 10610 10364 10674 10368
rect 10610 10308 10614 10364
rect 10614 10308 10670 10364
rect 10670 10308 10674 10364
rect 10610 10304 10674 10308
rect 2957 9820 3021 9824
rect 2957 9764 2961 9820
rect 2961 9764 3017 9820
rect 3017 9764 3021 9820
rect 2957 9760 3021 9764
rect 3037 9820 3101 9824
rect 3037 9764 3041 9820
rect 3041 9764 3097 9820
rect 3097 9764 3101 9820
rect 3037 9760 3101 9764
rect 3117 9820 3181 9824
rect 3117 9764 3121 9820
rect 3121 9764 3177 9820
rect 3177 9764 3181 9820
rect 3117 9760 3181 9764
rect 3197 9820 3261 9824
rect 3197 9764 3201 9820
rect 3201 9764 3257 9820
rect 3257 9764 3261 9820
rect 3197 9760 3261 9764
rect 5648 9820 5712 9824
rect 5648 9764 5652 9820
rect 5652 9764 5708 9820
rect 5708 9764 5712 9820
rect 5648 9760 5712 9764
rect 5728 9820 5792 9824
rect 5728 9764 5732 9820
rect 5732 9764 5788 9820
rect 5788 9764 5792 9820
rect 5728 9760 5792 9764
rect 5808 9820 5872 9824
rect 5808 9764 5812 9820
rect 5812 9764 5868 9820
rect 5868 9764 5872 9820
rect 5808 9760 5872 9764
rect 5888 9820 5952 9824
rect 5888 9764 5892 9820
rect 5892 9764 5948 9820
rect 5948 9764 5952 9820
rect 5888 9760 5952 9764
rect 8339 9820 8403 9824
rect 8339 9764 8343 9820
rect 8343 9764 8399 9820
rect 8399 9764 8403 9820
rect 8339 9760 8403 9764
rect 8419 9820 8483 9824
rect 8419 9764 8423 9820
rect 8423 9764 8479 9820
rect 8479 9764 8483 9820
rect 8419 9760 8483 9764
rect 8499 9820 8563 9824
rect 8499 9764 8503 9820
rect 8503 9764 8559 9820
rect 8559 9764 8563 9820
rect 8499 9760 8563 9764
rect 8579 9820 8643 9824
rect 8579 9764 8583 9820
rect 8583 9764 8639 9820
rect 8639 9764 8643 9820
rect 8579 9760 8643 9764
rect 11030 9820 11094 9824
rect 11030 9764 11034 9820
rect 11034 9764 11090 9820
rect 11090 9764 11094 9820
rect 11030 9760 11094 9764
rect 11110 9820 11174 9824
rect 11110 9764 11114 9820
rect 11114 9764 11170 9820
rect 11170 9764 11174 9820
rect 11110 9760 11174 9764
rect 11190 9820 11254 9824
rect 11190 9764 11194 9820
rect 11194 9764 11250 9820
rect 11250 9764 11254 9820
rect 11190 9760 11254 9764
rect 11270 9820 11334 9824
rect 11270 9764 11274 9820
rect 11274 9764 11330 9820
rect 11330 9764 11334 9820
rect 11270 9760 11334 9764
rect 2297 9276 2361 9280
rect 2297 9220 2301 9276
rect 2301 9220 2357 9276
rect 2357 9220 2361 9276
rect 2297 9216 2361 9220
rect 2377 9276 2441 9280
rect 2377 9220 2381 9276
rect 2381 9220 2437 9276
rect 2437 9220 2441 9276
rect 2377 9216 2441 9220
rect 2457 9276 2521 9280
rect 2457 9220 2461 9276
rect 2461 9220 2517 9276
rect 2517 9220 2521 9276
rect 2457 9216 2521 9220
rect 2537 9276 2601 9280
rect 2537 9220 2541 9276
rect 2541 9220 2597 9276
rect 2597 9220 2601 9276
rect 2537 9216 2601 9220
rect 4988 9276 5052 9280
rect 4988 9220 4992 9276
rect 4992 9220 5048 9276
rect 5048 9220 5052 9276
rect 4988 9216 5052 9220
rect 5068 9276 5132 9280
rect 5068 9220 5072 9276
rect 5072 9220 5128 9276
rect 5128 9220 5132 9276
rect 5068 9216 5132 9220
rect 5148 9276 5212 9280
rect 5148 9220 5152 9276
rect 5152 9220 5208 9276
rect 5208 9220 5212 9276
rect 5148 9216 5212 9220
rect 5228 9276 5292 9280
rect 5228 9220 5232 9276
rect 5232 9220 5288 9276
rect 5288 9220 5292 9276
rect 5228 9216 5292 9220
rect 7679 9276 7743 9280
rect 7679 9220 7683 9276
rect 7683 9220 7739 9276
rect 7739 9220 7743 9276
rect 7679 9216 7743 9220
rect 7759 9276 7823 9280
rect 7759 9220 7763 9276
rect 7763 9220 7819 9276
rect 7819 9220 7823 9276
rect 7759 9216 7823 9220
rect 7839 9276 7903 9280
rect 7839 9220 7843 9276
rect 7843 9220 7899 9276
rect 7899 9220 7903 9276
rect 7839 9216 7903 9220
rect 7919 9276 7983 9280
rect 7919 9220 7923 9276
rect 7923 9220 7979 9276
rect 7979 9220 7983 9276
rect 7919 9216 7983 9220
rect 10370 9276 10434 9280
rect 10370 9220 10374 9276
rect 10374 9220 10430 9276
rect 10430 9220 10434 9276
rect 10370 9216 10434 9220
rect 10450 9276 10514 9280
rect 10450 9220 10454 9276
rect 10454 9220 10510 9276
rect 10510 9220 10514 9276
rect 10450 9216 10514 9220
rect 10530 9276 10594 9280
rect 10530 9220 10534 9276
rect 10534 9220 10590 9276
rect 10590 9220 10594 9276
rect 10530 9216 10594 9220
rect 10610 9276 10674 9280
rect 10610 9220 10614 9276
rect 10614 9220 10670 9276
rect 10670 9220 10674 9276
rect 10610 9216 10674 9220
rect 2957 8732 3021 8736
rect 2957 8676 2961 8732
rect 2961 8676 3017 8732
rect 3017 8676 3021 8732
rect 2957 8672 3021 8676
rect 3037 8732 3101 8736
rect 3037 8676 3041 8732
rect 3041 8676 3097 8732
rect 3097 8676 3101 8732
rect 3037 8672 3101 8676
rect 3117 8732 3181 8736
rect 3117 8676 3121 8732
rect 3121 8676 3177 8732
rect 3177 8676 3181 8732
rect 3117 8672 3181 8676
rect 3197 8732 3261 8736
rect 3197 8676 3201 8732
rect 3201 8676 3257 8732
rect 3257 8676 3261 8732
rect 3197 8672 3261 8676
rect 5648 8732 5712 8736
rect 5648 8676 5652 8732
rect 5652 8676 5708 8732
rect 5708 8676 5712 8732
rect 5648 8672 5712 8676
rect 5728 8732 5792 8736
rect 5728 8676 5732 8732
rect 5732 8676 5788 8732
rect 5788 8676 5792 8732
rect 5728 8672 5792 8676
rect 5808 8732 5872 8736
rect 5808 8676 5812 8732
rect 5812 8676 5868 8732
rect 5868 8676 5872 8732
rect 5808 8672 5872 8676
rect 5888 8732 5952 8736
rect 5888 8676 5892 8732
rect 5892 8676 5948 8732
rect 5948 8676 5952 8732
rect 5888 8672 5952 8676
rect 8339 8732 8403 8736
rect 8339 8676 8343 8732
rect 8343 8676 8399 8732
rect 8399 8676 8403 8732
rect 8339 8672 8403 8676
rect 8419 8732 8483 8736
rect 8419 8676 8423 8732
rect 8423 8676 8479 8732
rect 8479 8676 8483 8732
rect 8419 8672 8483 8676
rect 8499 8732 8563 8736
rect 8499 8676 8503 8732
rect 8503 8676 8559 8732
rect 8559 8676 8563 8732
rect 8499 8672 8563 8676
rect 8579 8732 8643 8736
rect 8579 8676 8583 8732
rect 8583 8676 8639 8732
rect 8639 8676 8643 8732
rect 8579 8672 8643 8676
rect 11030 8732 11094 8736
rect 11030 8676 11034 8732
rect 11034 8676 11090 8732
rect 11090 8676 11094 8732
rect 11030 8672 11094 8676
rect 11110 8732 11174 8736
rect 11110 8676 11114 8732
rect 11114 8676 11170 8732
rect 11170 8676 11174 8732
rect 11110 8672 11174 8676
rect 11190 8732 11254 8736
rect 11190 8676 11194 8732
rect 11194 8676 11250 8732
rect 11250 8676 11254 8732
rect 11190 8672 11254 8676
rect 11270 8732 11334 8736
rect 11270 8676 11274 8732
rect 11274 8676 11330 8732
rect 11330 8676 11334 8732
rect 11270 8672 11334 8676
rect 2297 8188 2361 8192
rect 2297 8132 2301 8188
rect 2301 8132 2357 8188
rect 2357 8132 2361 8188
rect 2297 8128 2361 8132
rect 2377 8188 2441 8192
rect 2377 8132 2381 8188
rect 2381 8132 2437 8188
rect 2437 8132 2441 8188
rect 2377 8128 2441 8132
rect 2457 8188 2521 8192
rect 2457 8132 2461 8188
rect 2461 8132 2517 8188
rect 2517 8132 2521 8188
rect 2457 8128 2521 8132
rect 2537 8188 2601 8192
rect 2537 8132 2541 8188
rect 2541 8132 2597 8188
rect 2597 8132 2601 8188
rect 2537 8128 2601 8132
rect 4988 8188 5052 8192
rect 4988 8132 4992 8188
rect 4992 8132 5048 8188
rect 5048 8132 5052 8188
rect 4988 8128 5052 8132
rect 5068 8188 5132 8192
rect 5068 8132 5072 8188
rect 5072 8132 5128 8188
rect 5128 8132 5132 8188
rect 5068 8128 5132 8132
rect 5148 8188 5212 8192
rect 5148 8132 5152 8188
rect 5152 8132 5208 8188
rect 5208 8132 5212 8188
rect 5148 8128 5212 8132
rect 5228 8188 5292 8192
rect 5228 8132 5232 8188
rect 5232 8132 5288 8188
rect 5288 8132 5292 8188
rect 5228 8128 5292 8132
rect 7679 8188 7743 8192
rect 7679 8132 7683 8188
rect 7683 8132 7739 8188
rect 7739 8132 7743 8188
rect 7679 8128 7743 8132
rect 7759 8188 7823 8192
rect 7759 8132 7763 8188
rect 7763 8132 7819 8188
rect 7819 8132 7823 8188
rect 7759 8128 7823 8132
rect 7839 8188 7903 8192
rect 7839 8132 7843 8188
rect 7843 8132 7899 8188
rect 7899 8132 7903 8188
rect 7839 8128 7903 8132
rect 7919 8188 7983 8192
rect 7919 8132 7923 8188
rect 7923 8132 7979 8188
rect 7979 8132 7983 8188
rect 7919 8128 7983 8132
rect 10370 8188 10434 8192
rect 10370 8132 10374 8188
rect 10374 8132 10430 8188
rect 10430 8132 10434 8188
rect 10370 8128 10434 8132
rect 10450 8188 10514 8192
rect 10450 8132 10454 8188
rect 10454 8132 10510 8188
rect 10510 8132 10514 8188
rect 10450 8128 10514 8132
rect 10530 8188 10594 8192
rect 10530 8132 10534 8188
rect 10534 8132 10590 8188
rect 10590 8132 10594 8188
rect 10530 8128 10594 8132
rect 10610 8188 10674 8192
rect 10610 8132 10614 8188
rect 10614 8132 10670 8188
rect 10670 8132 10674 8188
rect 10610 8128 10674 8132
rect 2957 7644 3021 7648
rect 2957 7588 2961 7644
rect 2961 7588 3017 7644
rect 3017 7588 3021 7644
rect 2957 7584 3021 7588
rect 3037 7644 3101 7648
rect 3037 7588 3041 7644
rect 3041 7588 3097 7644
rect 3097 7588 3101 7644
rect 3037 7584 3101 7588
rect 3117 7644 3181 7648
rect 3117 7588 3121 7644
rect 3121 7588 3177 7644
rect 3177 7588 3181 7644
rect 3117 7584 3181 7588
rect 3197 7644 3261 7648
rect 3197 7588 3201 7644
rect 3201 7588 3257 7644
rect 3257 7588 3261 7644
rect 3197 7584 3261 7588
rect 5648 7644 5712 7648
rect 5648 7588 5652 7644
rect 5652 7588 5708 7644
rect 5708 7588 5712 7644
rect 5648 7584 5712 7588
rect 5728 7644 5792 7648
rect 5728 7588 5732 7644
rect 5732 7588 5788 7644
rect 5788 7588 5792 7644
rect 5728 7584 5792 7588
rect 5808 7644 5872 7648
rect 5808 7588 5812 7644
rect 5812 7588 5868 7644
rect 5868 7588 5872 7644
rect 5808 7584 5872 7588
rect 5888 7644 5952 7648
rect 5888 7588 5892 7644
rect 5892 7588 5948 7644
rect 5948 7588 5952 7644
rect 5888 7584 5952 7588
rect 8339 7644 8403 7648
rect 8339 7588 8343 7644
rect 8343 7588 8399 7644
rect 8399 7588 8403 7644
rect 8339 7584 8403 7588
rect 8419 7644 8483 7648
rect 8419 7588 8423 7644
rect 8423 7588 8479 7644
rect 8479 7588 8483 7644
rect 8419 7584 8483 7588
rect 8499 7644 8563 7648
rect 8499 7588 8503 7644
rect 8503 7588 8559 7644
rect 8559 7588 8563 7644
rect 8499 7584 8563 7588
rect 8579 7644 8643 7648
rect 8579 7588 8583 7644
rect 8583 7588 8639 7644
rect 8639 7588 8643 7644
rect 8579 7584 8643 7588
rect 11030 7644 11094 7648
rect 11030 7588 11034 7644
rect 11034 7588 11090 7644
rect 11090 7588 11094 7644
rect 11030 7584 11094 7588
rect 11110 7644 11174 7648
rect 11110 7588 11114 7644
rect 11114 7588 11170 7644
rect 11170 7588 11174 7644
rect 11110 7584 11174 7588
rect 11190 7644 11254 7648
rect 11190 7588 11194 7644
rect 11194 7588 11250 7644
rect 11250 7588 11254 7644
rect 11190 7584 11254 7588
rect 11270 7644 11334 7648
rect 11270 7588 11274 7644
rect 11274 7588 11330 7644
rect 11330 7588 11334 7644
rect 11270 7584 11334 7588
rect 2297 7100 2361 7104
rect 2297 7044 2301 7100
rect 2301 7044 2357 7100
rect 2357 7044 2361 7100
rect 2297 7040 2361 7044
rect 2377 7100 2441 7104
rect 2377 7044 2381 7100
rect 2381 7044 2437 7100
rect 2437 7044 2441 7100
rect 2377 7040 2441 7044
rect 2457 7100 2521 7104
rect 2457 7044 2461 7100
rect 2461 7044 2517 7100
rect 2517 7044 2521 7100
rect 2457 7040 2521 7044
rect 2537 7100 2601 7104
rect 2537 7044 2541 7100
rect 2541 7044 2597 7100
rect 2597 7044 2601 7100
rect 2537 7040 2601 7044
rect 4988 7100 5052 7104
rect 4988 7044 4992 7100
rect 4992 7044 5048 7100
rect 5048 7044 5052 7100
rect 4988 7040 5052 7044
rect 5068 7100 5132 7104
rect 5068 7044 5072 7100
rect 5072 7044 5128 7100
rect 5128 7044 5132 7100
rect 5068 7040 5132 7044
rect 5148 7100 5212 7104
rect 5148 7044 5152 7100
rect 5152 7044 5208 7100
rect 5208 7044 5212 7100
rect 5148 7040 5212 7044
rect 5228 7100 5292 7104
rect 5228 7044 5232 7100
rect 5232 7044 5288 7100
rect 5288 7044 5292 7100
rect 5228 7040 5292 7044
rect 7679 7100 7743 7104
rect 7679 7044 7683 7100
rect 7683 7044 7739 7100
rect 7739 7044 7743 7100
rect 7679 7040 7743 7044
rect 7759 7100 7823 7104
rect 7759 7044 7763 7100
rect 7763 7044 7819 7100
rect 7819 7044 7823 7100
rect 7759 7040 7823 7044
rect 7839 7100 7903 7104
rect 7839 7044 7843 7100
rect 7843 7044 7899 7100
rect 7899 7044 7903 7100
rect 7839 7040 7903 7044
rect 7919 7100 7983 7104
rect 7919 7044 7923 7100
rect 7923 7044 7979 7100
rect 7979 7044 7983 7100
rect 7919 7040 7983 7044
rect 10370 7100 10434 7104
rect 10370 7044 10374 7100
rect 10374 7044 10430 7100
rect 10430 7044 10434 7100
rect 10370 7040 10434 7044
rect 10450 7100 10514 7104
rect 10450 7044 10454 7100
rect 10454 7044 10510 7100
rect 10510 7044 10514 7100
rect 10450 7040 10514 7044
rect 10530 7100 10594 7104
rect 10530 7044 10534 7100
rect 10534 7044 10590 7100
rect 10590 7044 10594 7100
rect 10530 7040 10594 7044
rect 10610 7100 10674 7104
rect 10610 7044 10614 7100
rect 10614 7044 10670 7100
rect 10670 7044 10674 7100
rect 10610 7040 10674 7044
rect 6868 7032 6932 7036
rect 6868 6976 6918 7032
rect 6918 6976 6932 7032
rect 6868 6972 6932 6976
rect 9628 6972 9692 7036
rect 2957 6556 3021 6560
rect 2957 6500 2961 6556
rect 2961 6500 3017 6556
rect 3017 6500 3021 6556
rect 2957 6496 3021 6500
rect 3037 6556 3101 6560
rect 3037 6500 3041 6556
rect 3041 6500 3097 6556
rect 3097 6500 3101 6556
rect 3037 6496 3101 6500
rect 3117 6556 3181 6560
rect 3117 6500 3121 6556
rect 3121 6500 3177 6556
rect 3177 6500 3181 6556
rect 3117 6496 3181 6500
rect 3197 6556 3261 6560
rect 3197 6500 3201 6556
rect 3201 6500 3257 6556
rect 3257 6500 3261 6556
rect 3197 6496 3261 6500
rect 5648 6556 5712 6560
rect 5648 6500 5652 6556
rect 5652 6500 5708 6556
rect 5708 6500 5712 6556
rect 5648 6496 5712 6500
rect 5728 6556 5792 6560
rect 5728 6500 5732 6556
rect 5732 6500 5788 6556
rect 5788 6500 5792 6556
rect 5728 6496 5792 6500
rect 5808 6556 5872 6560
rect 5808 6500 5812 6556
rect 5812 6500 5868 6556
rect 5868 6500 5872 6556
rect 5808 6496 5872 6500
rect 5888 6556 5952 6560
rect 5888 6500 5892 6556
rect 5892 6500 5948 6556
rect 5948 6500 5952 6556
rect 5888 6496 5952 6500
rect 8339 6556 8403 6560
rect 8339 6500 8343 6556
rect 8343 6500 8399 6556
rect 8399 6500 8403 6556
rect 8339 6496 8403 6500
rect 8419 6556 8483 6560
rect 8419 6500 8423 6556
rect 8423 6500 8479 6556
rect 8479 6500 8483 6556
rect 8419 6496 8483 6500
rect 8499 6556 8563 6560
rect 8499 6500 8503 6556
rect 8503 6500 8559 6556
rect 8559 6500 8563 6556
rect 8499 6496 8563 6500
rect 8579 6556 8643 6560
rect 8579 6500 8583 6556
rect 8583 6500 8639 6556
rect 8639 6500 8643 6556
rect 8579 6496 8643 6500
rect 11030 6556 11094 6560
rect 11030 6500 11034 6556
rect 11034 6500 11090 6556
rect 11090 6500 11094 6556
rect 11030 6496 11094 6500
rect 11110 6556 11174 6560
rect 11110 6500 11114 6556
rect 11114 6500 11170 6556
rect 11170 6500 11174 6556
rect 11110 6496 11174 6500
rect 11190 6556 11254 6560
rect 11190 6500 11194 6556
rect 11194 6500 11250 6556
rect 11250 6500 11254 6556
rect 11190 6496 11254 6500
rect 11270 6556 11334 6560
rect 11270 6500 11274 6556
rect 11274 6500 11330 6556
rect 11330 6500 11334 6556
rect 11270 6496 11334 6500
rect 2297 6012 2361 6016
rect 2297 5956 2301 6012
rect 2301 5956 2357 6012
rect 2357 5956 2361 6012
rect 2297 5952 2361 5956
rect 2377 6012 2441 6016
rect 2377 5956 2381 6012
rect 2381 5956 2437 6012
rect 2437 5956 2441 6012
rect 2377 5952 2441 5956
rect 2457 6012 2521 6016
rect 2457 5956 2461 6012
rect 2461 5956 2517 6012
rect 2517 5956 2521 6012
rect 2457 5952 2521 5956
rect 2537 6012 2601 6016
rect 2537 5956 2541 6012
rect 2541 5956 2597 6012
rect 2597 5956 2601 6012
rect 2537 5952 2601 5956
rect 4988 6012 5052 6016
rect 4988 5956 4992 6012
rect 4992 5956 5048 6012
rect 5048 5956 5052 6012
rect 4988 5952 5052 5956
rect 5068 6012 5132 6016
rect 5068 5956 5072 6012
rect 5072 5956 5128 6012
rect 5128 5956 5132 6012
rect 5068 5952 5132 5956
rect 5148 6012 5212 6016
rect 5148 5956 5152 6012
rect 5152 5956 5208 6012
rect 5208 5956 5212 6012
rect 5148 5952 5212 5956
rect 5228 6012 5292 6016
rect 5228 5956 5232 6012
rect 5232 5956 5288 6012
rect 5288 5956 5292 6012
rect 5228 5952 5292 5956
rect 7679 6012 7743 6016
rect 7679 5956 7683 6012
rect 7683 5956 7739 6012
rect 7739 5956 7743 6012
rect 7679 5952 7743 5956
rect 7759 6012 7823 6016
rect 7759 5956 7763 6012
rect 7763 5956 7819 6012
rect 7819 5956 7823 6012
rect 7759 5952 7823 5956
rect 7839 6012 7903 6016
rect 7839 5956 7843 6012
rect 7843 5956 7899 6012
rect 7899 5956 7903 6012
rect 7839 5952 7903 5956
rect 7919 6012 7983 6016
rect 7919 5956 7923 6012
rect 7923 5956 7979 6012
rect 7979 5956 7983 6012
rect 7919 5952 7983 5956
rect 10370 6012 10434 6016
rect 10370 5956 10374 6012
rect 10374 5956 10430 6012
rect 10430 5956 10434 6012
rect 10370 5952 10434 5956
rect 10450 6012 10514 6016
rect 10450 5956 10454 6012
rect 10454 5956 10510 6012
rect 10510 5956 10514 6012
rect 10450 5952 10514 5956
rect 10530 6012 10594 6016
rect 10530 5956 10534 6012
rect 10534 5956 10590 6012
rect 10590 5956 10594 6012
rect 10530 5952 10594 5956
rect 10610 6012 10674 6016
rect 10610 5956 10614 6012
rect 10614 5956 10670 6012
rect 10670 5956 10674 6012
rect 10610 5952 10674 5956
rect 2957 5468 3021 5472
rect 2957 5412 2961 5468
rect 2961 5412 3017 5468
rect 3017 5412 3021 5468
rect 2957 5408 3021 5412
rect 3037 5468 3101 5472
rect 3037 5412 3041 5468
rect 3041 5412 3097 5468
rect 3097 5412 3101 5468
rect 3037 5408 3101 5412
rect 3117 5468 3181 5472
rect 3117 5412 3121 5468
rect 3121 5412 3177 5468
rect 3177 5412 3181 5468
rect 3117 5408 3181 5412
rect 3197 5468 3261 5472
rect 3197 5412 3201 5468
rect 3201 5412 3257 5468
rect 3257 5412 3261 5468
rect 3197 5408 3261 5412
rect 5648 5468 5712 5472
rect 5648 5412 5652 5468
rect 5652 5412 5708 5468
rect 5708 5412 5712 5468
rect 5648 5408 5712 5412
rect 5728 5468 5792 5472
rect 5728 5412 5732 5468
rect 5732 5412 5788 5468
rect 5788 5412 5792 5468
rect 5728 5408 5792 5412
rect 5808 5468 5872 5472
rect 5808 5412 5812 5468
rect 5812 5412 5868 5468
rect 5868 5412 5872 5468
rect 5808 5408 5872 5412
rect 5888 5468 5952 5472
rect 5888 5412 5892 5468
rect 5892 5412 5948 5468
rect 5948 5412 5952 5468
rect 5888 5408 5952 5412
rect 8339 5468 8403 5472
rect 8339 5412 8343 5468
rect 8343 5412 8399 5468
rect 8399 5412 8403 5468
rect 8339 5408 8403 5412
rect 8419 5468 8483 5472
rect 8419 5412 8423 5468
rect 8423 5412 8479 5468
rect 8479 5412 8483 5468
rect 8419 5408 8483 5412
rect 8499 5468 8563 5472
rect 8499 5412 8503 5468
rect 8503 5412 8559 5468
rect 8559 5412 8563 5468
rect 8499 5408 8563 5412
rect 8579 5468 8643 5472
rect 8579 5412 8583 5468
rect 8583 5412 8639 5468
rect 8639 5412 8643 5468
rect 8579 5408 8643 5412
rect 11030 5468 11094 5472
rect 11030 5412 11034 5468
rect 11034 5412 11090 5468
rect 11090 5412 11094 5468
rect 11030 5408 11094 5412
rect 11110 5468 11174 5472
rect 11110 5412 11114 5468
rect 11114 5412 11170 5468
rect 11170 5412 11174 5468
rect 11110 5408 11174 5412
rect 11190 5468 11254 5472
rect 11190 5412 11194 5468
rect 11194 5412 11250 5468
rect 11250 5412 11254 5468
rect 11190 5408 11254 5412
rect 11270 5468 11334 5472
rect 11270 5412 11274 5468
rect 11274 5412 11330 5468
rect 11330 5412 11334 5468
rect 11270 5408 11334 5412
rect 2297 4924 2361 4928
rect 2297 4868 2301 4924
rect 2301 4868 2357 4924
rect 2357 4868 2361 4924
rect 2297 4864 2361 4868
rect 2377 4924 2441 4928
rect 2377 4868 2381 4924
rect 2381 4868 2437 4924
rect 2437 4868 2441 4924
rect 2377 4864 2441 4868
rect 2457 4924 2521 4928
rect 2457 4868 2461 4924
rect 2461 4868 2517 4924
rect 2517 4868 2521 4924
rect 2457 4864 2521 4868
rect 2537 4924 2601 4928
rect 2537 4868 2541 4924
rect 2541 4868 2597 4924
rect 2597 4868 2601 4924
rect 2537 4864 2601 4868
rect 4988 4924 5052 4928
rect 4988 4868 4992 4924
rect 4992 4868 5048 4924
rect 5048 4868 5052 4924
rect 4988 4864 5052 4868
rect 5068 4924 5132 4928
rect 5068 4868 5072 4924
rect 5072 4868 5128 4924
rect 5128 4868 5132 4924
rect 5068 4864 5132 4868
rect 5148 4924 5212 4928
rect 5148 4868 5152 4924
rect 5152 4868 5208 4924
rect 5208 4868 5212 4924
rect 5148 4864 5212 4868
rect 5228 4924 5292 4928
rect 5228 4868 5232 4924
rect 5232 4868 5288 4924
rect 5288 4868 5292 4924
rect 5228 4864 5292 4868
rect 7679 4924 7743 4928
rect 7679 4868 7683 4924
rect 7683 4868 7739 4924
rect 7739 4868 7743 4924
rect 7679 4864 7743 4868
rect 7759 4924 7823 4928
rect 7759 4868 7763 4924
rect 7763 4868 7819 4924
rect 7819 4868 7823 4924
rect 7759 4864 7823 4868
rect 7839 4924 7903 4928
rect 7839 4868 7843 4924
rect 7843 4868 7899 4924
rect 7899 4868 7903 4924
rect 7839 4864 7903 4868
rect 7919 4924 7983 4928
rect 7919 4868 7923 4924
rect 7923 4868 7979 4924
rect 7979 4868 7983 4924
rect 7919 4864 7983 4868
rect 10370 4924 10434 4928
rect 10370 4868 10374 4924
rect 10374 4868 10430 4924
rect 10430 4868 10434 4924
rect 10370 4864 10434 4868
rect 10450 4924 10514 4928
rect 10450 4868 10454 4924
rect 10454 4868 10510 4924
rect 10510 4868 10514 4924
rect 10450 4864 10514 4868
rect 10530 4924 10594 4928
rect 10530 4868 10534 4924
rect 10534 4868 10590 4924
rect 10590 4868 10594 4924
rect 10530 4864 10594 4868
rect 10610 4924 10674 4928
rect 10610 4868 10614 4924
rect 10614 4868 10670 4924
rect 10670 4868 10674 4924
rect 10610 4864 10674 4868
rect 2957 4380 3021 4384
rect 2957 4324 2961 4380
rect 2961 4324 3017 4380
rect 3017 4324 3021 4380
rect 2957 4320 3021 4324
rect 3037 4380 3101 4384
rect 3037 4324 3041 4380
rect 3041 4324 3097 4380
rect 3097 4324 3101 4380
rect 3037 4320 3101 4324
rect 3117 4380 3181 4384
rect 3117 4324 3121 4380
rect 3121 4324 3177 4380
rect 3177 4324 3181 4380
rect 3117 4320 3181 4324
rect 3197 4380 3261 4384
rect 3197 4324 3201 4380
rect 3201 4324 3257 4380
rect 3257 4324 3261 4380
rect 3197 4320 3261 4324
rect 5648 4380 5712 4384
rect 5648 4324 5652 4380
rect 5652 4324 5708 4380
rect 5708 4324 5712 4380
rect 5648 4320 5712 4324
rect 5728 4380 5792 4384
rect 5728 4324 5732 4380
rect 5732 4324 5788 4380
rect 5788 4324 5792 4380
rect 5728 4320 5792 4324
rect 5808 4380 5872 4384
rect 5808 4324 5812 4380
rect 5812 4324 5868 4380
rect 5868 4324 5872 4380
rect 5808 4320 5872 4324
rect 5888 4380 5952 4384
rect 5888 4324 5892 4380
rect 5892 4324 5948 4380
rect 5948 4324 5952 4380
rect 5888 4320 5952 4324
rect 8339 4380 8403 4384
rect 8339 4324 8343 4380
rect 8343 4324 8399 4380
rect 8399 4324 8403 4380
rect 8339 4320 8403 4324
rect 8419 4380 8483 4384
rect 8419 4324 8423 4380
rect 8423 4324 8479 4380
rect 8479 4324 8483 4380
rect 8419 4320 8483 4324
rect 8499 4380 8563 4384
rect 8499 4324 8503 4380
rect 8503 4324 8559 4380
rect 8559 4324 8563 4380
rect 8499 4320 8563 4324
rect 8579 4380 8643 4384
rect 8579 4324 8583 4380
rect 8583 4324 8639 4380
rect 8639 4324 8643 4380
rect 8579 4320 8643 4324
rect 11030 4380 11094 4384
rect 11030 4324 11034 4380
rect 11034 4324 11090 4380
rect 11090 4324 11094 4380
rect 11030 4320 11094 4324
rect 11110 4380 11174 4384
rect 11110 4324 11114 4380
rect 11114 4324 11170 4380
rect 11170 4324 11174 4380
rect 11110 4320 11174 4324
rect 11190 4380 11254 4384
rect 11190 4324 11194 4380
rect 11194 4324 11250 4380
rect 11250 4324 11254 4380
rect 11190 4320 11254 4324
rect 11270 4380 11334 4384
rect 11270 4324 11274 4380
rect 11274 4324 11330 4380
rect 11330 4324 11334 4380
rect 11270 4320 11334 4324
rect 6868 3980 6932 4044
rect 2297 3836 2361 3840
rect 2297 3780 2301 3836
rect 2301 3780 2357 3836
rect 2357 3780 2361 3836
rect 2297 3776 2361 3780
rect 2377 3836 2441 3840
rect 2377 3780 2381 3836
rect 2381 3780 2437 3836
rect 2437 3780 2441 3836
rect 2377 3776 2441 3780
rect 2457 3836 2521 3840
rect 2457 3780 2461 3836
rect 2461 3780 2517 3836
rect 2517 3780 2521 3836
rect 2457 3776 2521 3780
rect 2537 3836 2601 3840
rect 2537 3780 2541 3836
rect 2541 3780 2597 3836
rect 2597 3780 2601 3836
rect 2537 3776 2601 3780
rect 4988 3836 5052 3840
rect 4988 3780 4992 3836
rect 4992 3780 5048 3836
rect 5048 3780 5052 3836
rect 4988 3776 5052 3780
rect 5068 3836 5132 3840
rect 5068 3780 5072 3836
rect 5072 3780 5128 3836
rect 5128 3780 5132 3836
rect 5068 3776 5132 3780
rect 5148 3836 5212 3840
rect 5148 3780 5152 3836
rect 5152 3780 5208 3836
rect 5208 3780 5212 3836
rect 5148 3776 5212 3780
rect 5228 3836 5292 3840
rect 5228 3780 5232 3836
rect 5232 3780 5288 3836
rect 5288 3780 5292 3836
rect 5228 3776 5292 3780
rect 7679 3836 7743 3840
rect 7679 3780 7683 3836
rect 7683 3780 7739 3836
rect 7739 3780 7743 3836
rect 7679 3776 7743 3780
rect 7759 3836 7823 3840
rect 7759 3780 7763 3836
rect 7763 3780 7819 3836
rect 7819 3780 7823 3836
rect 7759 3776 7823 3780
rect 7839 3836 7903 3840
rect 7839 3780 7843 3836
rect 7843 3780 7899 3836
rect 7899 3780 7903 3836
rect 7839 3776 7903 3780
rect 7919 3836 7983 3840
rect 7919 3780 7923 3836
rect 7923 3780 7979 3836
rect 7979 3780 7983 3836
rect 7919 3776 7983 3780
rect 10370 3836 10434 3840
rect 10370 3780 10374 3836
rect 10374 3780 10430 3836
rect 10430 3780 10434 3836
rect 10370 3776 10434 3780
rect 10450 3836 10514 3840
rect 10450 3780 10454 3836
rect 10454 3780 10510 3836
rect 10510 3780 10514 3836
rect 10450 3776 10514 3780
rect 10530 3836 10594 3840
rect 10530 3780 10534 3836
rect 10534 3780 10590 3836
rect 10590 3780 10594 3836
rect 10530 3776 10594 3780
rect 10610 3836 10674 3840
rect 10610 3780 10614 3836
rect 10614 3780 10670 3836
rect 10670 3780 10674 3836
rect 10610 3776 10674 3780
rect 9628 3436 9692 3500
rect 2957 3292 3021 3296
rect 2957 3236 2961 3292
rect 2961 3236 3017 3292
rect 3017 3236 3021 3292
rect 2957 3232 3021 3236
rect 3037 3292 3101 3296
rect 3037 3236 3041 3292
rect 3041 3236 3097 3292
rect 3097 3236 3101 3292
rect 3037 3232 3101 3236
rect 3117 3292 3181 3296
rect 3117 3236 3121 3292
rect 3121 3236 3177 3292
rect 3177 3236 3181 3292
rect 3117 3232 3181 3236
rect 3197 3292 3261 3296
rect 3197 3236 3201 3292
rect 3201 3236 3257 3292
rect 3257 3236 3261 3292
rect 3197 3232 3261 3236
rect 5648 3292 5712 3296
rect 5648 3236 5652 3292
rect 5652 3236 5708 3292
rect 5708 3236 5712 3292
rect 5648 3232 5712 3236
rect 5728 3292 5792 3296
rect 5728 3236 5732 3292
rect 5732 3236 5788 3292
rect 5788 3236 5792 3292
rect 5728 3232 5792 3236
rect 5808 3292 5872 3296
rect 5808 3236 5812 3292
rect 5812 3236 5868 3292
rect 5868 3236 5872 3292
rect 5808 3232 5872 3236
rect 5888 3292 5952 3296
rect 5888 3236 5892 3292
rect 5892 3236 5948 3292
rect 5948 3236 5952 3292
rect 5888 3232 5952 3236
rect 8339 3292 8403 3296
rect 8339 3236 8343 3292
rect 8343 3236 8399 3292
rect 8399 3236 8403 3292
rect 8339 3232 8403 3236
rect 8419 3292 8483 3296
rect 8419 3236 8423 3292
rect 8423 3236 8479 3292
rect 8479 3236 8483 3292
rect 8419 3232 8483 3236
rect 8499 3292 8563 3296
rect 8499 3236 8503 3292
rect 8503 3236 8559 3292
rect 8559 3236 8563 3292
rect 8499 3232 8563 3236
rect 8579 3292 8643 3296
rect 8579 3236 8583 3292
rect 8583 3236 8639 3292
rect 8639 3236 8643 3292
rect 8579 3232 8643 3236
rect 11030 3292 11094 3296
rect 11030 3236 11034 3292
rect 11034 3236 11090 3292
rect 11090 3236 11094 3292
rect 11030 3232 11094 3236
rect 11110 3292 11174 3296
rect 11110 3236 11114 3292
rect 11114 3236 11170 3292
rect 11170 3236 11174 3292
rect 11110 3232 11174 3236
rect 11190 3292 11254 3296
rect 11190 3236 11194 3292
rect 11194 3236 11250 3292
rect 11250 3236 11254 3292
rect 11190 3232 11254 3236
rect 11270 3292 11334 3296
rect 11270 3236 11274 3292
rect 11274 3236 11330 3292
rect 11330 3236 11334 3292
rect 11270 3232 11334 3236
rect 2297 2748 2361 2752
rect 2297 2692 2301 2748
rect 2301 2692 2357 2748
rect 2357 2692 2361 2748
rect 2297 2688 2361 2692
rect 2377 2748 2441 2752
rect 2377 2692 2381 2748
rect 2381 2692 2437 2748
rect 2437 2692 2441 2748
rect 2377 2688 2441 2692
rect 2457 2748 2521 2752
rect 2457 2692 2461 2748
rect 2461 2692 2517 2748
rect 2517 2692 2521 2748
rect 2457 2688 2521 2692
rect 2537 2748 2601 2752
rect 2537 2692 2541 2748
rect 2541 2692 2597 2748
rect 2597 2692 2601 2748
rect 2537 2688 2601 2692
rect 4988 2748 5052 2752
rect 4988 2692 4992 2748
rect 4992 2692 5048 2748
rect 5048 2692 5052 2748
rect 4988 2688 5052 2692
rect 5068 2748 5132 2752
rect 5068 2692 5072 2748
rect 5072 2692 5128 2748
rect 5128 2692 5132 2748
rect 5068 2688 5132 2692
rect 5148 2748 5212 2752
rect 5148 2692 5152 2748
rect 5152 2692 5208 2748
rect 5208 2692 5212 2748
rect 5148 2688 5212 2692
rect 5228 2748 5292 2752
rect 5228 2692 5232 2748
rect 5232 2692 5288 2748
rect 5288 2692 5292 2748
rect 5228 2688 5292 2692
rect 7679 2748 7743 2752
rect 7679 2692 7683 2748
rect 7683 2692 7739 2748
rect 7739 2692 7743 2748
rect 7679 2688 7743 2692
rect 7759 2748 7823 2752
rect 7759 2692 7763 2748
rect 7763 2692 7819 2748
rect 7819 2692 7823 2748
rect 7759 2688 7823 2692
rect 7839 2748 7903 2752
rect 7839 2692 7843 2748
rect 7843 2692 7899 2748
rect 7899 2692 7903 2748
rect 7839 2688 7903 2692
rect 7919 2748 7983 2752
rect 7919 2692 7923 2748
rect 7923 2692 7979 2748
rect 7979 2692 7983 2748
rect 7919 2688 7983 2692
rect 10370 2748 10434 2752
rect 10370 2692 10374 2748
rect 10374 2692 10430 2748
rect 10430 2692 10434 2748
rect 10370 2688 10434 2692
rect 10450 2748 10514 2752
rect 10450 2692 10454 2748
rect 10454 2692 10510 2748
rect 10510 2692 10514 2748
rect 10450 2688 10514 2692
rect 10530 2748 10594 2752
rect 10530 2692 10534 2748
rect 10534 2692 10590 2748
rect 10590 2692 10594 2748
rect 10530 2688 10594 2692
rect 10610 2748 10674 2752
rect 10610 2692 10614 2748
rect 10614 2692 10670 2748
rect 10670 2692 10674 2748
rect 10610 2688 10674 2692
rect 2957 2204 3021 2208
rect 2957 2148 2961 2204
rect 2961 2148 3017 2204
rect 3017 2148 3021 2204
rect 2957 2144 3021 2148
rect 3037 2204 3101 2208
rect 3037 2148 3041 2204
rect 3041 2148 3097 2204
rect 3097 2148 3101 2204
rect 3037 2144 3101 2148
rect 3117 2204 3181 2208
rect 3117 2148 3121 2204
rect 3121 2148 3177 2204
rect 3177 2148 3181 2204
rect 3117 2144 3181 2148
rect 3197 2204 3261 2208
rect 3197 2148 3201 2204
rect 3201 2148 3257 2204
rect 3257 2148 3261 2204
rect 3197 2144 3261 2148
rect 5648 2204 5712 2208
rect 5648 2148 5652 2204
rect 5652 2148 5708 2204
rect 5708 2148 5712 2204
rect 5648 2144 5712 2148
rect 5728 2204 5792 2208
rect 5728 2148 5732 2204
rect 5732 2148 5788 2204
rect 5788 2148 5792 2204
rect 5728 2144 5792 2148
rect 5808 2204 5872 2208
rect 5808 2148 5812 2204
rect 5812 2148 5868 2204
rect 5868 2148 5872 2204
rect 5808 2144 5872 2148
rect 5888 2204 5952 2208
rect 5888 2148 5892 2204
rect 5892 2148 5948 2204
rect 5948 2148 5952 2204
rect 5888 2144 5952 2148
rect 8339 2204 8403 2208
rect 8339 2148 8343 2204
rect 8343 2148 8399 2204
rect 8399 2148 8403 2204
rect 8339 2144 8403 2148
rect 8419 2204 8483 2208
rect 8419 2148 8423 2204
rect 8423 2148 8479 2204
rect 8479 2148 8483 2204
rect 8419 2144 8483 2148
rect 8499 2204 8563 2208
rect 8499 2148 8503 2204
rect 8503 2148 8559 2204
rect 8559 2148 8563 2204
rect 8499 2144 8563 2148
rect 8579 2204 8643 2208
rect 8579 2148 8583 2204
rect 8583 2148 8639 2204
rect 8639 2148 8643 2204
rect 8579 2144 8643 2148
rect 11030 2204 11094 2208
rect 11030 2148 11034 2204
rect 11034 2148 11090 2204
rect 11090 2148 11094 2204
rect 11030 2144 11094 2148
rect 11110 2204 11174 2208
rect 11110 2148 11114 2204
rect 11114 2148 11170 2204
rect 11170 2148 11174 2204
rect 11110 2144 11174 2148
rect 11190 2204 11254 2208
rect 11190 2148 11194 2204
rect 11194 2148 11250 2204
rect 11250 2148 11254 2204
rect 11190 2144 11254 2148
rect 11270 2204 11334 2208
rect 11270 2148 11274 2204
rect 11274 2148 11330 2204
rect 11330 2148 11334 2204
rect 11270 2144 11334 2148
<< metal4 >>
rect 2289 12544 2609 12560
rect 2289 12480 2297 12544
rect 2361 12480 2377 12544
rect 2441 12480 2457 12544
rect 2521 12480 2537 12544
rect 2601 12480 2609 12544
rect 2289 11456 2609 12480
rect 2289 11392 2297 11456
rect 2361 11392 2377 11456
rect 2441 11392 2457 11456
rect 2521 11392 2537 11456
rect 2601 11392 2609 11456
rect 2289 11338 2609 11392
rect 2289 11102 2331 11338
rect 2567 11102 2609 11338
rect 2289 10368 2609 11102
rect 2289 10304 2297 10368
rect 2361 10304 2377 10368
rect 2441 10304 2457 10368
rect 2521 10304 2537 10368
rect 2601 10304 2609 10368
rect 2289 9280 2609 10304
rect 2289 9216 2297 9280
rect 2361 9216 2377 9280
rect 2441 9216 2457 9280
rect 2521 9216 2537 9280
rect 2601 9216 2609 9280
rect 2289 8754 2609 9216
rect 2289 8518 2331 8754
rect 2567 8518 2609 8754
rect 2289 8192 2609 8518
rect 2289 8128 2297 8192
rect 2361 8128 2377 8192
rect 2441 8128 2457 8192
rect 2521 8128 2537 8192
rect 2601 8128 2609 8192
rect 2289 7104 2609 8128
rect 2289 7040 2297 7104
rect 2361 7040 2377 7104
rect 2441 7040 2457 7104
rect 2521 7040 2537 7104
rect 2601 7040 2609 7104
rect 2289 6170 2609 7040
rect 2289 6016 2331 6170
rect 2567 6016 2609 6170
rect 2289 5952 2297 6016
rect 2601 5952 2609 6016
rect 2289 5934 2331 5952
rect 2567 5934 2609 5952
rect 2289 4928 2609 5934
rect 2289 4864 2297 4928
rect 2361 4864 2377 4928
rect 2441 4864 2457 4928
rect 2521 4864 2537 4928
rect 2601 4864 2609 4928
rect 2289 3840 2609 4864
rect 2289 3776 2297 3840
rect 2361 3776 2377 3840
rect 2441 3776 2457 3840
rect 2521 3776 2537 3840
rect 2601 3776 2609 3840
rect 2289 3586 2609 3776
rect 2289 3350 2331 3586
rect 2567 3350 2609 3586
rect 2289 2752 2609 3350
rect 2289 2688 2297 2752
rect 2361 2688 2377 2752
rect 2441 2688 2457 2752
rect 2521 2688 2537 2752
rect 2601 2688 2609 2752
rect 2289 2128 2609 2688
rect 2949 12000 3269 12560
rect 2949 11936 2957 12000
rect 3021 11998 3037 12000
rect 3101 11998 3117 12000
rect 3181 11998 3197 12000
rect 3261 11936 3269 12000
rect 2949 11762 2991 11936
rect 3227 11762 3269 11936
rect 2949 10912 3269 11762
rect 2949 10848 2957 10912
rect 3021 10848 3037 10912
rect 3101 10848 3117 10912
rect 3181 10848 3197 10912
rect 3261 10848 3269 10912
rect 2949 9824 3269 10848
rect 2949 9760 2957 9824
rect 3021 9760 3037 9824
rect 3101 9760 3117 9824
rect 3181 9760 3197 9824
rect 3261 9760 3269 9824
rect 2949 9414 3269 9760
rect 2949 9178 2991 9414
rect 3227 9178 3269 9414
rect 2949 8736 3269 9178
rect 2949 8672 2957 8736
rect 3021 8672 3037 8736
rect 3101 8672 3117 8736
rect 3181 8672 3197 8736
rect 3261 8672 3269 8736
rect 2949 7648 3269 8672
rect 2949 7584 2957 7648
rect 3021 7584 3037 7648
rect 3101 7584 3117 7648
rect 3181 7584 3197 7648
rect 3261 7584 3269 7648
rect 2949 6830 3269 7584
rect 2949 6594 2991 6830
rect 3227 6594 3269 6830
rect 2949 6560 3269 6594
rect 2949 6496 2957 6560
rect 3021 6496 3037 6560
rect 3101 6496 3117 6560
rect 3181 6496 3197 6560
rect 3261 6496 3269 6560
rect 2949 5472 3269 6496
rect 2949 5408 2957 5472
rect 3021 5408 3037 5472
rect 3101 5408 3117 5472
rect 3181 5408 3197 5472
rect 3261 5408 3269 5472
rect 2949 4384 3269 5408
rect 2949 4320 2957 4384
rect 3021 4320 3037 4384
rect 3101 4320 3117 4384
rect 3181 4320 3197 4384
rect 3261 4320 3269 4384
rect 2949 4246 3269 4320
rect 2949 4010 2991 4246
rect 3227 4010 3269 4246
rect 2949 3296 3269 4010
rect 2949 3232 2957 3296
rect 3021 3232 3037 3296
rect 3101 3232 3117 3296
rect 3181 3232 3197 3296
rect 3261 3232 3269 3296
rect 2949 2208 3269 3232
rect 2949 2144 2957 2208
rect 3021 2144 3037 2208
rect 3101 2144 3117 2208
rect 3181 2144 3197 2208
rect 3261 2144 3269 2208
rect 2949 2128 3269 2144
rect 4980 12544 5300 12560
rect 4980 12480 4988 12544
rect 5052 12480 5068 12544
rect 5132 12480 5148 12544
rect 5212 12480 5228 12544
rect 5292 12480 5300 12544
rect 4980 11456 5300 12480
rect 4980 11392 4988 11456
rect 5052 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5300 11456
rect 4980 11338 5300 11392
rect 4980 11102 5022 11338
rect 5258 11102 5300 11338
rect 4980 10368 5300 11102
rect 4980 10304 4988 10368
rect 5052 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5300 10368
rect 4980 9280 5300 10304
rect 4980 9216 4988 9280
rect 5052 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5300 9280
rect 4980 8754 5300 9216
rect 4980 8518 5022 8754
rect 5258 8518 5300 8754
rect 4980 8192 5300 8518
rect 4980 8128 4988 8192
rect 5052 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5300 8192
rect 4980 7104 5300 8128
rect 4980 7040 4988 7104
rect 5052 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5300 7104
rect 4980 6170 5300 7040
rect 4980 6016 5022 6170
rect 5258 6016 5300 6170
rect 4980 5952 4988 6016
rect 5292 5952 5300 6016
rect 4980 5934 5022 5952
rect 5258 5934 5300 5952
rect 4980 4928 5300 5934
rect 4980 4864 4988 4928
rect 5052 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5300 4928
rect 4980 3840 5300 4864
rect 4980 3776 4988 3840
rect 5052 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5300 3840
rect 4980 3586 5300 3776
rect 4980 3350 5022 3586
rect 5258 3350 5300 3586
rect 4980 2752 5300 3350
rect 4980 2688 4988 2752
rect 5052 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5300 2752
rect 4980 2128 5300 2688
rect 5640 12000 5960 12560
rect 5640 11936 5648 12000
rect 5712 11998 5728 12000
rect 5792 11998 5808 12000
rect 5872 11998 5888 12000
rect 5952 11936 5960 12000
rect 5640 11762 5682 11936
rect 5918 11762 5960 11936
rect 5640 10912 5960 11762
rect 5640 10848 5648 10912
rect 5712 10848 5728 10912
rect 5792 10848 5808 10912
rect 5872 10848 5888 10912
rect 5952 10848 5960 10912
rect 5640 9824 5960 10848
rect 5640 9760 5648 9824
rect 5712 9760 5728 9824
rect 5792 9760 5808 9824
rect 5872 9760 5888 9824
rect 5952 9760 5960 9824
rect 5640 9414 5960 9760
rect 5640 9178 5682 9414
rect 5918 9178 5960 9414
rect 5640 8736 5960 9178
rect 5640 8672 5648 8736
rect 5712 8672 5728 8736
rect 5792 8672 5808 8736
rect 5872 8672 5888 8736
rect 5952 8672 5960 8736
rect 5640 7648 5960 8672
rect 5640 7584 5648 7648
rect 5712 7584 5728 7648
rect 5792 7584 5808 7648
rect 5872 7584 5888 7648
rect 5952 7584 5960 7648
rect 5640 6830 5960 7584
rect 7671 12544 7991 12560
rect 7671 12480 7679 12544
rect 7743 12480 7759 12544
rect 7823 12480 7839 12544
rect 7903 12480 7919 12544
rect 7983 12480 7991 12544
rect 7671 11456 7991 12480
rect 7671 11392 7679 11456
rect 7743 11392 7759 11456
rect 7823 11392 7839 11456
rect 7903 11392 7919 11456
rect 7983 11392 7991 11456
rect 7671 11338 7991 11392
rect 7671 11102 7713 11338
rect 7949 11102 7991 11338
rect 7671 10368 7991 11102
rect 7671 10304 7679 10368
rect 7743 10304 7759 10368
rect 7823 10304 7839 10368
rect 7903 10304 7919 10368
rect 7983 10304 7991 10368
rect 7671 9280 7991 10304
rect 7671 9216 7679 9280
rect 7743 9216 7759 9280
rect 7823 9216 7839 9280
rect 7903 9216 7919 9280
rect 7983 9216 7991 9280
rect 7671 8754 7991 9216
rect 7671 8518 7713 8754
rect 7949 8518 7991 8754
rect 7671 8192 7991 8518
rect 7671 8128 7679 8192
rect 7743 8128 7759 8192
rect 7823 8128 7839 8192
rect 7903 8128 7919 8192
rect 7983 8128 7991 8192
rect 7671 7104 7991 8128
rect 7671 7040 7679 7104
rect 7743 7040 7759 7104
rect 7823 7040 7839 7104
rect 7903 7040 7919 7104
rect 7983 7040 7991 7104
rect 6867 7036 6933 7037
rect 6867 6972 6868 7036
rect 6932 6972 6933 7036
rect 6867 6971 6933 6972
rect 5640 6594 5682 6830
rect 5918 6594 5960 6830
rect 5640 6560 5960 6594
rect 5640 6496 5648 6560
rect 5712 6496 5728 6560
rect 5792 6496 5808 6560
rect 5872 6496 5888 6560
rect 5952 6496 5960 6560
rect 5640 5472 5960 6496
rect 5640 5408 5648 5472
rect 5712 5408 5728 5472
rect 5792 5408 5808 5472
rect 5872 5408 5888 5472
rect 5952 5408 5960 5472
rect 5640 4384 5960 5408
rect 5640 4320 5648 4384
rect 5712 4320 5728 4384
rect 5792 4320 5808 4384
rect 5872 4320 5888 4384
rect 5952 4320 5960 4384
rect 5640 4246 5960 4320
rect 5640 4010 5682 4246
rect 5918 4010 5960 4246
rect 6870 4045 6930 6971
rect 7671 6170 7991 7040
rect 7671 6016 7713 6170
rect 7949 6016 7991 6170
rect 7671 5952 7679 6016
rect 7983 5952 7991 6016
rect 7671 5934 7713 5952
rect 7949 5934 7991 5952
rect 7671 4928 7991 5934
rect 7671 4864 7679 4928
rect 7743 4864 7759 4928
rect 7823 4864 7839 4928
rect 7903 4864 7919 4928
rect 7983 4864 7991 4928
rect 5640 3296 5960 4010
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 5640 3232 5648 3296
rect 5712 3232 5728 3296
rect 5792 3232 5808 3296
rect 5872 3232 5888 3296
rect 5952 3232 5960 3296
rect 5640 2208 5960 3232
rect 5640 2144 5648 2208
rect 5712 2144 5728 2208
rect 5792 2144 5808 2208
rect 5872 2144 5888 2208
rect 5952 2144 5960 2208
rect 5640 2128 5960 2144
rect 7671 3840 7991 4864
rect 7671 3776 7679 3840
rect 7743 3776 7759 3840
rect 7823 3776 7839 3840
rect 7903 3776 7919 3840
rect 7983 3776 7991 3840
rect 7671 3586 7991 3776
rect 7671 3350 7713 3586
rect 7949 3350 7991 3586
rect 7671 2752 7991 3350
rect 7671 2688 7679 2752
rect 7743 2688 7759 2752
rect 7823 2688 7839 2752
rect 7903 2688 7919 2752
rect 7983 2688 7991 2752
rect 7671 2128 7991 2688
rect 8331 12000 8651 12560
rect 8331 11936 8339 12000
rect 8403 11998 8419 12000
rect 8483 11998 8499 12000
rect 8563 11998 8579 12000
rect 8643 11936 8651 12000
rect 8331 11762 8373 11936
rect 8609 11762 8651 11936
rect 8331 10912 8651 11762
rect 8331 10848 8339 10912
rect 8403 10848 8419 10912
rect 8483 10848 8499 10912
rect 8563 10848 8579 10912
rect 8643 10848 8651 10912
rect 8331 9824 8651 10848
rect 8331 9760 8339 9824
rect 8403 9760 8419 9824
rect 8483 9760 8499 9824
rect 8563 9760 8579 9824
rect 8643 9760 8651 9824
rect 8331 9414 8651 9760
rect 8331 9178 8373 9414
rect 8609 9178 8651 9414
rect 8331 8736 8651 9178
rect 8331 8672 8339 8736
rect 8403 8672 8419 8736
rect 8483 8672 8499 8736
rect 8563 8672 8579 8736
rect 8643 8672 8651 8736
rect 8331 7648 8651 8672
rect 8331 7584 8339 7648
rect 8403 7584 8419 7648
rect 8483 7584 8499 7648
rect 8563 7584 8579 7648
rect 8643 7584 8651 7648
rect 8331 6830 8651 7584
rect 10362 12544 10682 12560
rect 10362 12480 10370 12544
rect 10434 12480 10450 12544
rect 10514 12480 10530 12544
rect 10594 12480 10610 12544
rect 10674 12480 10682 12544
rect 10362 11456 10682 12480
rect 10362 11392 10370 11456
rect 10434 11392 10450 11456
rect 10514 11392 10530 11456
rect 10594 11392 10610 11456
rect 10674 11392 10682 11456
rect 10362 11338 10682 11392
rect 10362 11102 10404 11338
rect 10640 11102 10682 11338
rect 10362 10368 10682 11102
rect 10362 10304 10370 10368
rect 10434 10304 10450 10368
rect 10514 10304 10530 10368
rect 10594 10304 10610 10368
rect 10674 10304 10682 10368
rect 10362 9280 10682 10304
rect 10362 9216 10370 9280
rect 10434 9216 10450 9280
rect 10514 9216 10530 9280
rect 10594 9216 10610 9280
rect 10674 9216 10682 9280
rect 10362 8754 10682 9216
rect 10362 8518 10404 8754
rect 10640 8518 10682 8754
rect 10362 8192 10682 8518
rect 10362 8128 10370 8192
rect 10434 8128 10450 8192
rect 10514 8128 10530 8192
rect 10594 8128 10610 8192
rect 10674 8128 10682 8192
rect 10362 7104 10682 8128
rect 10362 7040 10370 7104
rect 10434 7040 10450 7104
rect 10514 7040 10530 7104
rect 10594 7040 10610 7104
rect 10674 7040 10682 7104
rect 9627 7036 9693 7037
rect 9627 6972 9628 7036
rect 9692 6972 9693 7036
rect 9627 6971 9693 6972
rect 8331 6594 8373 6830
rect 8609 6594 8651 6830
rect 8331 6560 8651 6594
rect 8331 6496 8339 6560
rect 8403 6496 8419 6560
rect 8483 6496 8499 6560
rect 8563 6496 8579 6560
rect 8643 6496 8651 6560
rect 8331 5472 8651 6496
rect 8331 5408 8339 5472
rect 8403 5408 8419 5472
rect 8483 5408 8499 5472
rect 8563 5408 8579 5472
rect 8643 5408 8651 5472
rect 8331 4384 8651 5408
rect 8331 4320 8339 4384
rect 8403 4320 8419 4384
rect 8483 4320 8499 4384
rect 8563 4320 8579 4384
rect 8643 4320 8651 4384
rect 8331 4246 8651 4320
rect 8331 4010 8373 4246
rect 8609 4010 8651 4246
rect 8331 3296 8651 4010
rect 9630 3501 9690 6971
rect 10362 6170 10682 7040
rect 10362 6016 10404 6170
rect 10640 6016 10682 6170
rect 10362 5952 10370 6016
rect 10674 5952 10682 6016
rect 10362 5934 10404 5952
rect 10640 5934 10682 5952
rect 10362 4928 10682 5934
rect 10362 4864 10370 4928
rect 10434 4864 10450 4928
rect 10514 4864 10530 4928
rect 10594 4864 10610 4928
rect 10674 4864 10682 4928
rect 10362 3840 10682 4864
rect 10362 3776 10370 3840
rect 10434 3776 10450 3840
rect 10514 3776 10530 3840
rect 10594 3776 10610 3840
rect 10674 3776 10682 3840
rect 10362 3586 10682 3776
rect 9627 3500 9693 3501
rect 9627 3436 9628 3500
rect 9692 3436 9693 3500
rect 9627 3435 9693 3436
rect 8331 3232 8339 3296
rect 8403 3232 8419 3296
rect 8483 3232 8499 3296
rect 8563 3232 8579 3296
rect 8643 3232 8651 3296
rect 8331 2208 8651 3232
rect 8331 2144 8339 2208
rect 8403 2144 8419 2208
rect 8483 2144 8499 2208
rect 8563 2144 8579 2208
rect 8643 2144 8651 2208
rect 8331 2128 8651 2144
rect 10362 3350 10404 3586
rect 10640 3350 10682 3586
rect 10362 2752 10682 3350
rect 10362 2688 10370 2752
rect 10434 2688 10450 2752
rect 10514 2688 10530 2752
rect 10594 2688 10610 2752
rect 10674 2688 10682 2752
rect 10362 2128 10682 2688
rect 11022 12000 11342 12560
rect 11022 11936 11030 12000
rect 11094 11998 11110 12000
rect 11174 11998 11190 12000
rect 11254 11998 11270 12000
rect 11334 11936 11342 12000
rect 11022 11762 11064 11936
rect 11300 11762 11342 11936
rect 11022 10912 11342 11762
rect 11022 10848 11030 10912
rect 11094 10848 11110 10912
rect 11174 10848 11190 10912
rect 11254 10848 11270 10912
rect 11334 10848 11342 10912
rect 11022 9824 11342 10848
rect 11022 9760 11030 9824
rect 11094 9760 11110 9824
rect 11174 9760 11190 9824
rect 11254 9760 11270 9824
rect 11334 9760 11342 9824
rect 11022 9414 11342 9760
rect 11022 9178 11064 9414
rect 11300 9178 11342 9414
rect 11022 8736 11342 9178
rect 11022 8672 11030 8736
rect 11094 8672 11110 8736
rect 11174 8672 11190 8736
rect 11254 8672 11270 8736
rect 11334 8672 11342 8736
rect 11022 7648 11342 8672
rect 11022 7584 11030 7648
rect 11094 7584 11110 7648
rect 11174 7584 11190 7648
rect 11254 7584 11270 7648
rect 11334 7584 11342 7648
rect 11022 6830 11342 7584
rect 11022 6594 11064 6830
rect 11300 6594 11342 6830
rect 11022 6560 11342 6594
rect 11022 6496 11030 6560
rect 11094 6496 11110 6560
rect 11174 6496 11190 6560
rect 11254 6496 11270 6560
rect 11334 6496 11342 6560
rect 11022 5472 11342 6496
rect 11022 5408 11030 5472
rect 11094 5408 11110 5472
rect 11174 5408 11190 5472
rect 11254 5408 11270 5472
rect 11334 5408 11342 5472
rect 11022 4384 11342 5408
rect 11022 4320 11030 4384
rect 11094 4320 11110 4384
rect 11174 4320 11190 4384
rect 11254 4320 11270 4384
rect 11334 4320 11342 4384
rect 11022 4246 11342 4320
rect 11022 4010 11064 4246
rect 11300 4010 11342 4246
rect 11022 3296 11342 4010
rect 11022 3232 11030 3296
rect 11094 3232 11110 3296
rect 11174 3232 11190 3296
rect 11254 3232 11270 3296
rect 11334 3232 11342 3296
rect 11022 2208 11342 3232
rect 11022 2144 11030 2208
rect 11094 2144 11110 2208
rect 11174 2144 11190 2208
rect 11254 2144 11270 2208
rect 11334 2144 11342 2208
rect 11022 2128 11342 2144
<< via4 >>
rect 2331 11102 2567 11338
rect 2331 8518 2567 8754
rect 2331 6016 2567 6170
rect 2331 5952 2361 6016
rect 2361 5952 2377 6016
rect 2377 5952 2441 6016
rect 2441 5952 2457 6016
rect 2457 5952 2521 6016
rect 2521 5952 2537 6016
rect 2537 5952 2567 6016
rect 2331 5934 2567 5952
rect 2331 3350 2567 3586
rect 2991 11936 3021 11998
rect 3021 11936 3037 11998
rect 3037 11936 3101 11998
rect 3101 11936 3117 11998
rect 3117 11936 3181 11998
rect 3181 11936 3197 11998
rect 3197 11936 3227 11998
rect 2991 11762 3227 11936
rect 2991 9178 3227 9414
rect 2991 6594 3227 6830
rect 2991 4010 3227 4246
rect 5022 11102 5258 11338
rect 5022 8518 5258 8754
rect 5022 6016 5258 6170
rect 5022 5952 5052 6016
rect 5052 5952 5068 6016
rect 5068 5952 5132 6016
rect 5132 5952 5148 6016
rect 5148 5952 5212 6016
rect 5212 5952 5228 6016
rect 5228 5952 5258 6016
rect 5022 5934 5258 5952
rect 5022 3350 5258 3586
rect 5682 11936 5712 11998
rect 5712 11936 5728 11998
rect 5728 11936 5792 11998
rect 5792 11936 5808 11998
rect 5808 11936 5872 11998
rect 5872 11936 5888 11998
rect 5888 11936 5918 11998
rect 5682 11762 5918 11936
rect 5682 9178 5918 9414
rect 7713 11102 7949 11338
rect 7713 8518 7949 8754
rect 5682 6594 5918 6830
rect 5682 4010 5918 4246
rect 7713 6016 7949 6170
rect 7713 5952 7743 6016
rect 7743 5952 7759 6016
rect 7759 5952 7823 6016
rect 7823 5952 7839 6016
rect 7839 5952 7903 6016
rect 7903 5952 7919 6016
rect 7919 5952 7949 6016
rect 7713 5934 7949 5952
rect 7713 3350 7949 3586
rect 8373 11936 8403 11998
rect 8403 11936 8419 11998
rect 8419 11936 8483 11998
rect 8483 11936 8499 11998
rect 8499 11936 8563 11998
rect 8563 11936 8579 11998
rect 8579 11936 8609 11998
rect 8373 11762 8609 11936
rect 8373 9178 8609 9414
rect 10404 11102 10640 11338
rect 10404 8518 10640 8754
rect 8373 6594 8609 6830
rect 8373 4010 8609 4246
rect 10404 6016 10640 6170
rect 10404 5952 10434 6016
rect 10434 5952 10450 6016
rect 10450 5952 10514 6016
rect 10514 5952 10530 6016
rect 10530 5952 10594 6016
rect 10594 5952 10610 6016
rect 10610 5952 10640 6016
rect 10404 5934 10640 5952
rect 10404 3350 10640 3586
rect 11064 11936 11094 11998
rect 11094 11936 11110 11998
rect 11110 11936 11174 11998
rect 11174 11936 11190 11998
rect 11190 11936 11254 11998
rect 11254 11936 11270 11998
rect 11270 11936 11300 11998
rect 11064 11762 11300 11936
rect 11064 9178 11300 9414
rect 11064 6594 11300 6830
rect 11064 4010 11300 4246
<< metal5 >>
rect 1056 11998 11916 12040
rect 1056 11762 2991 11998
rect 3227 11762 5682 11998
rect 5918 11762 8373 11998
rect 8609 11762 11064 11998
rect 11300 11762 11916 11998
rect 1056 11720 11916 11762
rect 1056 11338 11916 11380
rect 1056 11102 2331 11338
rect 2567 11102 5022 11338
rect 5258 11102 7713 11338
rect 7949 11102 10404 11338
rect 10640 11102 11916 11338
rect 1056 11060 11916 11102
rect 1056 9414 11916 9456
rect 1056 9178 2991 9414
rect 3227 9178 5682 9414
rect 5918 9178 8373 9414
rect 8609 9178 11064 9414
rect 11300 9178 11916 9414
rect 1056 9136 11916 9178
rect 1056 8754 11916 8796
rect 1056 8518 2331 8754
rect 2567 8518 5022 8754
rect 5258 8518 7713 8754
rect 7949 8518 10404 8754
rect 10640 8518 11916 8754
rect 1056 8476 11916 8518
rect 1056 6830 11916 6872
rect 1056 6594 2991 6830
rect 3227 6594 5682 6830
rect 5918 6594 8373 6830
rect 8609 6594 11064 6830
rect 11300 6594 11916 6830
rect 1056 6552 11916 6594
rect 1056 6170 11916 6212
rect 1056 5934 2331 6170
rect 2567 5934 5022 6170
rect 5258 5934 7713 6170
rect 7949 5934 10404 6170
rect 10640 5934 11916 6170
rect 1056 5892 11916 5934
rect 1056 4246 11916 4288
rect 1056 4010 2991 4246
rect 3227 4010 5682 4246
rect 5918 4010 8373 4246
rect 8609 4010 11064 4246
rect 11300 4010 11916 4246
rect 1056 3968 11916 4010
rect 1056 3586 11916 3628
rect 1056 3350 2331 3586
rect 2567 3350 5022 3586
rect 5258 3350 7713 3586
rect 7949 3350 10404 3586
rect 10640 3350 11916 3586
rect 1056 3308 11916 3350
use sky130_fd_sc_hd__clkbuf_4  _121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _122_
timestamp 1723858470
transform 1 0 4140 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _123_
timestamp 1723858470
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7636 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _126_
timestamp 1723858470
transform -1 0 6716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9568 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _130_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9292 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _131_
timestamp 1723858470
transform -1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _132_
timestamp 1723858470
transform 1 0 3864 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 2668 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _134_
timestamp 1723858470
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _135_
timestamp 1723858470
transform -1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _136_
timestamp 1723858470
transform 1 0 2392 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _137_
timestamp 1723858470
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _138_
timestamp 1723858470
transform 1 0 2392 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _139_
timestamp 1723858470
transform -1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 3404 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_2  _142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1748 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _144_
timestamp 1723858470
transform 1 0 1564 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _145_
timestamp 1723858470
transform -1 0 3496 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _146_
timestamp 1723858470
transform -1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _147_
timestamp 1723858470
transform -1 0 3680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2944 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o41ai_1  _150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5888 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _151_
timestamp 1723858470
transform -1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _152_
timestamp 1723858470
transform 1 0 6716 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _153_
timestamp 1723858470
transform -1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6900 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _156_
timestamp 1723858470
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _157_
timestamp 1723858470
transform 1 0 8372 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9384 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8832 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _161_
timestamp 1723858470
transform -1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_2  _162_
timestamp 1723858470
transform 1 0 8924 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _164_
timestamp 1723858470
transform 1 0 4876 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _165_
timestamp 1723858470
transform 1 0 5428 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _166_
timestamp 1723858470
transform 1 0 4692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5428 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5520 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1723858470
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _170_
timestamp 1723858470
transform 1 0 7820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _171_
timestamp 1723858470
transform 1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _174_
timestamp 1723858470
transform 1 0 8832 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _175_
timestamp 1723858470
transform -1 0 10396 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1723858470
transform 1 0 10396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _177_
timestamp 1723858470
transform 1 0 8648 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _178_
timestamp 1723858470
transform -1 0 10304 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1723858470
transform 1 0 9936 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _180_
timestamp 1723858470
transform -1 0 8372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _181_
timestamp 1723858470
transform -1 0 8740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _182_
timestamp 1723858470
transform 1 0 9384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9384 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _184_
timestamp 1723858470
transform -1 0 10212 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1723858470
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1723858470
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _188_
timestamp 1723858470
transform 1 0 9016 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9660 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _190_
timestamp 1723858470
transform 1 0 6440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _191_
timestamp 1723858470
transform -1 0 8188 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _192_
timestamp 1723858470
transform 1 0 6900 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1723858470
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _194_
timestamp 1723858470
transform -1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7544 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _196_
timestamp 1723858470
transform 1 0 6348 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _197_
timestamp 1723858470
transform -1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _198_
timestamp 1723858470
transform -1 0 5612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _199_
timestamp 1723858470
transform -1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _200_
timestamp 1723858470
transform 1 0 3036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _201_
timestamp 1723858470
transform 1 0 1932 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _202_
timestamp 1723858470
transform 1 0 1932 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1723858470
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _204_
timestamp 1723858470
transform 1 0 3496 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 1723858470
transform -1 0 5152 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1723858470
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4416 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _208_
timestamp 1723858470
transform 1 0 3496 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1723858470
transform -1 0 4968 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1723858470
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _211_
timestamp 1723858470
transform 1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _212_
timestamp 1723858470
transform -1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _213_
timestamp 1723858470
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _214_
timestamp 1723858470
transform 1 0 2852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _215_
timestamp 1723858470
transform 1 0 1840 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1723858470
transform -1 0 2760 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1723858470
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1723858470
transform 1 0 3312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _219_
timestamp 1723858470
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3404 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _221_
timestamp 1723858470
transform 1 0 4048 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _222_
timestamp 1723858470
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _223_
timestamp 1723858470
transform 1 0 2116 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _224_
timestamp 1723858470
transform 1 0 8188 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1723858470
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1723858470
transform -1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1723858470
transform -1 0 4784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1723858470
transform -1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1723858470
transform -1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1723858470
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1723858470
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1723858470
transform -1 0 3680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1723858470
transform 1 0 6900 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1723858470
transform 1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1723858470
transform -1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1723858470
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1723858470
transform -1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1723858470
transform -1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1723858470
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1723858470
transform -1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8832 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 3220 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _244_
timestamp 1723858470
transform -1 0 4876 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1656 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _246_
timestamp 1723858470
transform 1 0 4140 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _247_
timestamp 1723858470
transform -1 0 6072 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _248_
timestamp 1723858470
transform 1 0 4876 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _249_
timestamp 1723858470
transform 1 0 1564 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _250_
timestamp 1723858470
transform 1 0 6348 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _251_
timestamp 1723858470
transform 1 0 6256 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _252_
timestamp 1723858470
transform 1 0 9476 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _253_
timestamp 1723858470
transform 1 0 7728 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _254_
timestamp 1723858470
transform 1 0 9568 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _255_
timestamp 1723858470
transform 1 0 9568 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _256_
timestamp 1723858470
transform 1 0 6716 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _257_
timestamp 1723858470
transform 1 0 4876 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8188 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1723858470
transform -1 0 6256 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1723858470
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 1723858470
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1723858470
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_70 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1723858470
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_91
timestamp 1723858470
transform 1 0 9476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_103 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 1723858470
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_3
timestamp 1723858470
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_32
timestamp 1723858470
transform 1 0 4048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 1723858470
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_92
timestamp 1723858470
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_104
timestamp 1723858470
transform 1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1723858470
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_21
timestamp 1723858470
transform 1 0 3036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_29
timestamp 1723858470
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_35
timestamp 1723858470
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_77
timestamp 1723858470
transform 1 0 8188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1723858470
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_94
timestamp 1723858470
transform 1 0 9752 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 1723858470
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_25
timestamp 1723858470
transform 1 0 3404 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1723858470
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1723858470
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1723858470
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1723858470
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_81
timestamp 1723858470
transform 1 0 8556 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_86
timestamp 1723858470
transform 1 0 9016 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_98
timestamp 1723858470
transform 1 0 10120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1723858470
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1723858470
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_3
timestamp 1723858470
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_12
timestamp 1723858470
transform 1 0 2208 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_24
timestamp 1723858470
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_29
timestamp 1723858470
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_35
timestamp 1723858470
transform 1 0 4324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_42
timestamp 1723858470
transform 1 0 4968 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_48
timestamp 1723858470
transform 1 0 5520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_57
timestamp 1723858470
transform 1 0 6348 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1723858470
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1723858470
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_99
timestamp 1723858470
transform 1 0 10212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_111
timestamp 1723858470
transform 1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 1723858470
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_30
timestamp 1723858470
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_36
timestamp 1723858470
transform 1 0 4416 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_40
timestamp 1723858470
transform 1 0 4784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1723858470
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_63
timestamp 1723858470
transform 1 0 6900 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_75
timestamp 1723858470
transform 1 0 8004 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_94
timestamp 1723858470
transform 1 0 9752 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_106
timestamp 1723858470
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1723858470
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1723858470
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_20
timestamp 1723858470
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1723858470
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_49
timestamp 1723858470
transform 1 0 5612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_61
timestamp 1723858470
transform 1 0 6716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_73
timestamp 1723858470
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_98
timestamp 1723858470
transform 1 0 10120 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_104
timestamp 1723858470
transform 1 0 10672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_3
timestamp 1723858470
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_16
timestamp 1723858470
transform 1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_27
timestamp 1723858470
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_34
timestamp 1723858470
transform 1 0 4232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_52
timestamp 1723858470
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 1723858470
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_72
timestamp 1723858470
transform 1 0 7728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1723858470
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1723858470
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_12
timestamp 1723858470
transform 1 0 2208 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_20
timestamp 1723858470
transform 1 0 2944 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1723858470
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_41
timestamp 1723858470
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_49
timestamp 1723858470
transform 1 0 5612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_73
timestamp 1723858470
transform 1 0 7820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_79
timestamp 1723858470
transform 1 0 8372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1723858470
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_100
timestamp 1723858470
transform 1 0 10304 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_112
timestamp 1723858470
transform 1 0 11408 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1723858470
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_15
timestamp 1723858470
transform 1 0 2484 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1723858470
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1723858470
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1723858470
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_77
timestamp 1723858470
transform 1 0 8188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_89
timestamp 1723858470
transform 1 0 9292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_101
timestamp 1723858470
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 1723858470
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1723858470
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1723858470
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_17
timestamp 1723858470
transform 1 0 2668 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1723858470
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_41
timestamp 1723858470
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_65
timestamp 1723858470
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_69
timestamp 1723858470
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_104
timestamp 1723858470
transform 1 0 10672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_108
timestamp 1723858470
transform 1 0 11040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1723858470
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_7
timestamp 1723858470
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_15
timestamp 1723858470
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_24
timestamp 1723858470
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_30
timestamp 1723858470
transform 1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_34
timestamp 1723858470
transform 1 0 4232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_47
timestamp 1723858470
transform 1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_51
timestamp 1723858470
transform 1 0 5796 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1723858470
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_78
timestamp 1723858470
transform 1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_91
timestamp 1723858470
transform 1 0 9476 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1723858470
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_6
timestamp 1723858470
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_15
timestamp 1723858470
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_39
timestamp 1723858470
transform 1 0 4692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_62
timestamp 1723858470
transform 1 0 6808 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_66
timestamp 1723858470
transform 1 0 7176 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_102
timestamp 1723858470
transform 1 0 10488 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1723858470
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_11
timestamp 1723858470
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_19
timestamp 1723858470
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_31
timestamp 1723858470
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_43
timestamp 1723858470
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1723858470
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1723858470
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1723858470
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_81
timestamp 1723858470
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_97
timestamp 1723858470
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1723858470
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1723858470
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 1723858470
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_11
timestamp 1723858470
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_22
timestamp 1723858470
transform 1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1723858470
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_35
timestamp 1723858470
transform 1 0 4324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_44
timestamp 1723858470
transform 1 0 5152 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_54
timestamp 1723858470
transform 1 0 6072 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 1723858470
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1723858470
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_85
timestamp 1723858470
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_100
timestamp 1723858470
transform 1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_104
timestamp 1723858470
transform 1 0 10672 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1723858470
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_11
timestamp 1723858470
transform 1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_45
timestamp 1723858470
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1723858470
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_82
timestamp 1723858470
transform 1 0 8648 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_90
timestamp 1723858470
transform 1 0 9384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 1723858470
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1723858470
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_40
timestamp 1723858470
transform 1 0 4784 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_99
timestamp 1723858470
transform 1 0 10212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_111
timestamp 1723858470
transform 1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_9
timestamp 1723858470
transform 1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_19
timestamp 1723858470
transform 1 0 2852 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1723858470
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1723858470
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1723858470
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_62
timestamp 1723858470
transform 1 0 6808 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_74
timestamp 1723858470
transform 1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_105
timestamp 1723858470
transform 1 0 10764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_113
timestamp 1723858470
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_7
timestamp 1723858470
transform 1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_25
timestamp 1723858470
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1723858470
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1723858470
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_44
timestamp 1723858470
transform 1 0 5152 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_57
timestamp 1723858470
transform 1 0 6348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_69
timestamp 1723858470
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_79
timestamp 1723858470
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1723858470
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_85
timestamp 1723858470
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_91
timestamp 1723858470
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_100
timestamp 1723858470
transform 1 0 10304 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_107
timestamp 1723858470
transform 1 0 10948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_113
timestamp 1723858470
transform 1 0 11500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 10304 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1723858470
transform -1 0 9660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1723858470
transform 1 0 2116 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1723858470
transform -1 0 8280 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1723858470
transform -1 0 4508 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1723858470
transform -1 0 6348 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1723858470
transform -1 0 11592 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1723858470
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1723858470
transform -1 0 8372 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1723858470
transform -1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1723858470
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1723858470
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1723858470
transform -1 0 1932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1723858470
transform -1 0 5152 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1723858470
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1723858470
transform -1 0 3404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1723858470
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1723858470
transform -1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1723858470
transform -1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1723858470
transform 1 0 11040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1723858470
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1723858470
transform 1 0 10396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1723858470
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1723858470
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1723858470
transform -1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1723858470
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1723858470
transform -1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1723858470
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1723858470
transform -1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1723858470
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1723858470
transform -1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1723858470
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1723858470
transform -1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1723858470
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1723858470
transform -1 0 11868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1723858470
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1723858470
transform -1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1723858470
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1723858470
transform -1 0 11868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1723858470
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1723858470
transform -1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1723858470
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1723858470
transform -1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1723858470
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1723858470
transform -1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1723858470
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1723858470
transform -1 0 11868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1723858470
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1723858470
transform -1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1723858470
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1723858470
transform -1 0 11868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1723858470
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1723858470
transform -1 0 11868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1723858470
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1723858470
transform -1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1723858470
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1723858470
transform -1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1723858470
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1723858470
transform -1 0 11868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1723858470
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1723858470
transform -1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1723858470
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1723858470
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1723858470
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1723858470
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1723858470
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1723858470
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1723858470
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1723858470
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1723858470
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1723858470
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1723858470
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1723858470
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1723858470
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1723858470
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1723858470
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1723858470
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1723858470
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1723858470
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1723858470
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1723858470
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1723858470
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1723858470
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1723858470
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1723858470
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1723858470
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1723858470
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1723858470
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1723858470
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1723858470
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1723858470
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1723858470
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1723858470
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1723858470
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1723858470
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1723858470
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1723858470
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1723858470
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1723858470
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1723858470
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1723858470
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1723858470
transform 1 0 11408 0 1 11968
box -38 -48 130 592
<< labels >>
flabel metal4 s 2949 2128 3269 12560 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5640 2128 5960 12560 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8331 2128 8651 12560 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11022 2128 11342 12560 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3968 11916 4288 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6552 11916 6872 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9136 11916 9456 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 11720 11916 12040 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2289 2128 2609 12560 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4980 2128 5300 12560 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7671 2128 7991 12560 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10362 2128 10682 12560 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3308 11916 3628 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5892 11916 6212 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8476 11916 8796 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 11060 11916 11380 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 12202 3408 13002 3528 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 12898 14346 12954 15146 0 FreeSans 224 90 0 0 count[0]
port 3 nsew signal tristate
flabel metal2 s 7746 14346 7802 15146 0 FreeSans 224 90 0 0 count[10]
port 4 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 count[11]
port 5 nsew signal tristate
flabel metal3 s 12202 12248 13002 12368 0 FreeSans 480 0 0 0 count[12]
port 6 nsew signal tristate
flabel metal3 s 12202 688 13002 808 0 FreeSans 480 0 0 0 count[13]
port 7 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 count[14]
port 8 nsew signal tristate
flabel metal2 s 4526 14346 4582 15146 0 FreeSans 224 90 0 0 count[15]
port 9 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 count[1]
port 10 nsew signal tristate
flabel metal2 s 1950 14346 2006 15146 0 FreeSans 224 90 0 0 count[2]
port 11 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 count[3]
port 12 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 count[4]
port 13 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 count[5]
port 14 nsew signal tristate
flabel metal3 s 12202 9528 13002 9648 0 FreeSans 480 0 0 0 count[6]
port 15 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 count[7]
port 16 nsew signal tristate
flabel metal2 s 10322 14346 10378 15146 0 FreeSans 224 90 0 0 count[8]
port 17 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 count[9]
port 18 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 ctrl
port 19 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 en
port 20 nsew signal input
flabel metal3 s 12202 6128 13002 6248 0 FreeSans 480 0 0 0 rst
port 21 nsew signal input
rlabel metal1 6486 11968 6486 11968 0 VGND
rlabel metal1 6486 12512 6486 12512 0 VPWR
rlabel metal2 9798 11560 9798 11560 0 _000_
rlabel metal2 2438 10914 2438 10914 0 _001_
rlabel metal1 4370 11322 4370 11322 0 _002_
rlabel metal1 3549 3094 3549 3094 0 _003_
rlabel metal1 5428 3910 5428 3910 0 _004_
rlabel metal1 5343 2346 5343 2346 0 _005_
rlabel metal1 6118 8602 6118 8602 0 _006_
rlabel metal2 3542 3944 3542 3944 0 _007_
rlabel metal2 7130 8670 7130 8670 0 _008_
rlabel metal1 7360 2618 7360 2618 0 _009_
rlabel metal2 10902 6086 10902 6086 0 _010_
rlabel metal2 8786 3502 8786 3502 0 _011_
rlabel metal2 10902 10472 10902 10472 0 _012_
rlabel metal2 10902 8296 10902 8296 0 _013_
rlabel metal1 8471 11050 8471 11050 0 _014_
rlabel metal1 6493 11118 6493 11118 0 _015_
rlabel metal1 8786 11730 8786 11730 0 _016_
rlabel metal2 2162 11356 2162 11356 0 _017_
rlabel metal1 4278 10778 4278 10778 0 _018_
rlabel metal2 2714 3026 2714 3026 0 _019_
rlabel metal1 4508 3094 4508 3094 0 _020_
rlabel metal2 5750 2621 5750 2621 0 _021_
rlabel metal2 5198 8738 5198 8738 0 _022_
rlabel metal1 1932 4182 1932 4182 0 _023_
rlabel metal1 6486 6630 6486 6630 0 _024_
rlabel metal1 6624 3162 6624 3162 0 _025_
rlabel metal1 9798 6392 9798 6392 0 _026_
rlabel metal1 8096 2958 8096 2958 0 _027_
rlabel metal1 9936 10710 9936 10710 0 _028_
rlabel metal1 10350 8058 10350 8058 0 _029_
rlabel metal1 7084 10778 7084 10778 0 _030_
rlabel metal1 5421 11322 5421 11322 0 _031_
rlabel metal2 5106 5780 5106 5780 0 _032_
rlabel metal1 7314 10540 7314 10540 0 _033_
rlabel metal1 7544 10234 7544 10234 0 _034_
rlabel metal1 8970 8466 8970 8466 0 _035_
rlabel metal2 9890 8092 9890 8092 0 _036_
rlabel metal1 10488 7854 10488 7854 0 _037_
rlabel metal1 9476 9486 9476 9486 0 _038_
rlabel metal1 10212 10234 10212 10234 0 _039_
rlabel metal2 8970 6154 8970 6154 0 _040_
rlabel metal1 8970 5712 8970 5712 0 _041_
rlabel metal1 9522 5746 9522 5746 0 _042_
rlabel metal2 10074 5100 10074 5100 0 _043_
rlabel metal1 9522 3502 9522 3502 0 _044_
rlabel metal1 8786 3502 8786 3502 0 _045_
rlabel metal1 9614 5882 9614 5882 0 _046_
rlabel metal1 9476 6426 9476 6426 0 _047_
rlabel metal1 7498 4658 7498 4658 0 _048_
rlabel metal1 7498 3162 7498 3162 0 _049_
rlabel metal1 6900 3026 6900 3026 0 _050_
rlabel metal1 7084 6834 7084 6834 0 _051_
rlabel metal1 6762 6766 6762 6766 0 _052_
rlabel metal1 4554 5168 4554 5168 0 _053_
rlabel metal1 4968 5542 4968 5542 0 _054_
rlabel metal1 3358 6800 3358 6800 0 _055_
rlabel metal1 2254 6324 2254 6324 0 _056_
rlabel metal1 2576 5338 2576 5338 0 _057_
rlabel metal1 2070 4590 2070 4590 0 _058_
rlabel metal1 4370 7310 4370 7310 0 _059_
rlabel metal1 5244 8466 5244 8466 0 _060_
rlabel metal2 3818 4250 3818 4250 0 _061_
rlabel metal1 4278 3978 4278 3978 0 _062_
rlabel metal1 4968 4114 4968 4114 0 _063_
rlabel metal2 4738 5508 4738 5508 0 _064_
rlabel metal2 4830 5882 4830 5882 0 _065_
rlabel metal1 2898 8500 2898 8500 0 _066_
rlabel metal1 2208 3502 2208 3502 0 _067_
rlabel metal1 2714 3434 2714 3434 0 _068_
rlabel metal1 3542 10234 3542 10234 0 _069_
rlabel metal1 3680 10166 3680 10166 0 _070_
rlabel metal1 3634 10506 3634 10506 0 _071_
rlabel metal1 2438 11662 2438 11662 0 _072_
rlabel via2 2530 10659 2530 10659 0 _073_
rlabel metal1 1932 5746 1932 5746 0 _074_
rlabel metal2 8694 7072 8694 7072 0 _075_
rlabel metal1 7406 9996 7406 9996 0 _076_
rlabel metal1 6808 10642 6808 10642 0 _077_
rlabel metal1 6670 10676 6670 10676 0 _078_
rlabel metal1 6762 10778 6762 10778 0 _079_
rlabel metal2 9062 8262 9062 8262 0 _080_
rlabel metal1 8786 8534 8786 8534 0 _081_
rlabel metal1 10258 8874 10258 8874 0 _082_
rlabel metal1 10442 9010 10442 9010 0 _083_
rlabel metal1 9338 8976 9338 8976 0 _084_
rlabel metal1 4646 6256 4646 6256 0 _085_
rlabel metal1 1932 8466 1932 8466 0 _086_
rlabel metal1 3312 8330 3312 8330 0 _087_
rlabel metal1 3082 8908 3082 8908 0 _088_
rlabel metal1 3496 8942 3496 8942 0 _089_
rlabel metal1 3542 10064 3542 10064 0 _090_
rlabel metal1 3358 11118 3358 11118 0 _091_
rlabel metal1 3220 10642 3220 10642 0 _092_
rlabel metal1 3726 9146 3726 9146 0 _093_
rlabel metal1 4232 8602 4232 8602 0 _094_
rlabel metal1 4830 6324 4830 6324 0 _095_
rlabel metal1 3312 5542 3312 5542 0 _096_
rlabel metal1 2162 6188 2162 6188 0 _097_
rlabel metal1 3266 7514 3266 7514 0 _098_
rlabel metal2 3634 7412 3634 7412 0 _099_
rlabel metal1 3634 7378 3634 7378 0 _100_
rlabel metal1 4922 6392 4922 6392 0 _101_
rlabel metal1 5842 6698 5842 6698 0 _102_
rlabel metal1 6440 6426 6440 6426 0 _103_
rlabel metal1 7314 6188 7314 6188 0 _104_
rlabel metal1 7682 6324 7682 6324 0 _105_
rlabel metal1 6808 6698 6808 6698 0 _106_
rlabel metal1 6486 6324 6486 6324 0 _107_
rlabel metal1 8878 5202 8878 5202 0 _108_
rlabel metal1 9338 4794 9338 4794 0 _109_
rlabel metal2 9062 5916 9062 5916 0 _110_
rlabel metal1 8970 5338 8970 5338 0 _111_
rlabel metal1 9016 5814 9016 5814 0 _112_
rlabel metal2 9430 7786 9430 7786 0 _113_
rlabel metal1 9844 8874 9844 8874 0 _114_
rlabel metal1 9568 9078 9568 9078 0 _115_
rlabel metal1 6210 10030 6210 10030 0 _116_
rlabel metal2 5474 11305 5474 11305 0 _117_
rlabel metal2 5934 10404 5934 10404 0 _118_
rlabel metal1 7636 2958 7636 2958 0 _119_
rlabel metal1 5428 10778 5428 10778 0 _120_
rlabel metal1 8188 7378 8188 7378 0 clk
rlabel metal1 6900 7174 6900 7174 0 clknet_0_clk
rlabel metal1 7314 3570 7314 3570 0 clknet_1_0__leaf_clk
rlabel metal2 9614 9520 9614 9520 0 clknet_1_1__leaf_clk
rlabel metal1 12098 11866 12098 11866 0 count[0]
rlabel metal2 7919 14484 7919 14484 0 count[10]
rlabel metal2 5198 823 5198 823 0 count[11]
rlabel metal2 11270 12359 11270 12359 0 count[12]
rlabel metal1 10994 2278 10994 2278 0 count[13]
rlabel metal3 820 11628 820 11628 0 count[14]
rlabel metal2 4554 13445 4554 13445 0 count[15]
rlabel metal2 46 1554 46 1554 0 count[1]
rlabel metal2 1978 13440 1978 13440 0 count[2]
rlabel metal2 10994 1112 10994 1112 0 count[3]
rlabel metal2 2622 1520 2622 1520 0 count[4]
rlabel metal3 820 2788 820 2788 0 count[5]
rlabel metal1 11776 9894 11776 9894 0 count[6]
rlabel metal3 820 5508 820 5508 0 count[7]
rlabel metal2 10297 14484 10297 14484 0 count[8]
rlabel metal2 8418 823 8418 823 0 count[9]
rlabel metal3 820 8908 820 8908 0 ctrl
rlabel metal3 843 14348 843 14348 0 en
rlabel metal2 2070 8364 2070 8364 0 net1
rlabel metal1 5060 11730 5060 11730 0 net10
rlabel metal1 1840 2414 1840 2414 0 net11
rlabel metal1 3082 8500 3082 8500 0 net12
rlabel metal2 2346 3094 2346 3094 0 net13
rlabel metal1 3726 2414 3726 2414 0 net14
rlabel metal2 2714 3944 2714 3944 0 net15
rlabel metal1 7774 9146 7774 9146 0 net16
rlabel metal1 3496 5270 3496 5270 0 net17
rlabel metal1 8188 12070 8188 12070 0 net18
rlabel metal1 8648 2414 8648 2414 0 net19
rlabel metal1 2300 5134 2300 5134 0 net2
rlabel metal1 8602 11662 8602 11662 0 net20
rlabel metal1 8372 10710 8372 10710 0 net21
rlabel metal1 2806 11798 2806 11798 0 net22
rlabel metal1 7176 6766 7176 6766 0 net23
rlabel metal2 3818 10812 3818 10812 0 net24
rlabel metal1 5612 4794 5612 4794 0 net25
rlabel metal1 8556 11118 8556 11118 0 net3
rlabel metal1 10396 11866 10396 11866 0 net4
rlabel metal1 8464 6290 8464 6290 0 net5
rlabel metal1 8142 2346 8142 2346 0 net6
rlabel metal1 11408 10778 11408 10778 0 net7
rlabel metal1 10902 2414 10902 2414 0 net8
rlabel metal1 2024 11798 2024 11798 0 net9
rlabel metal1 11638 5678 11638 5678 0 rst
<< properties >>
string FIXED_BBOX 0 0 13002 15146
<< end >>
