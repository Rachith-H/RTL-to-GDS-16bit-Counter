* NGSPICE file created from counter_up_dwn.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

.subckt counter_up_dwn VGND VPWR clk count[0] count[10] count[11] count[12] count[13]
+ count[14] count[15] count[1] count[2] count[3] count[4] count[5] count[6] count[7]
+ count[8] count[9] ctrl en rst
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_200_ _100_ _055_ _098_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__a21oi_1
X_131_ _082_ _083_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput7 net7 VGND VGND VPWR VPWR count[12] sky130_fd_sc_hd__buf_2
XFILLER_0_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_130_ net7 _076_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput10 net10 VGND VGND VPWR VPWR count[15] sky130_fd_sc_hd__clkbuf_4
Xoutput8 net8 VGND VGND VPWR VPWR count[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_189_ _119_ _042_ _046_ _047_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput11 net11 VGND VGND VPWR VPWR count[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR count[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_188_ _032_ net5 VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__and2_1
X_257_ clknet_1_1__leaf_clk _031_ _015_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
Xoutput12 net12 VGND VGND VPWR VPWR count[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_187_ _110_ _040_ _041_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__or3_1
X_256_ clknet_1_1__leaf_clk _030_ _014_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_239_ net3 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput13 net13 VGND VGND VPWR VPWR count[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_186_ _045_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__clkbuf_1
X_255_ clknet_1_1__leaf_clk _029_ _013_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfrtp_1
X_169_ net2 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__inv_2
X_238_ net3 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__inv_2
Xoutput14 net14 VGND VGND VPWR VPWR count[4] sky130_fd_sc_hd__clkbuf_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_185_ net6 _044_ _119_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__mux2_1
X_254_ clknet_1_1__leaf_clk _028_ _012_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_168_ _120_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__clkbuf_1
X_237_ net3 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__inv_2
Xoutput15 net15 VGND VGND VPWR VPWR count[5] sky130_fd_sc_hd__clkbuf_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_253_ clknet_1_0__leaf_clk _027_ _011_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfrtp_1
X_184_ _109_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__xnor2_1
X_236_ net3 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
X_167_ net10 _118_ _119_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ _090_ _093_ _119_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__o21a_1
Xoutput16 net16 VGND VGND VPWR VPWR count[6] sky130_fd_sc_hd__clkbuf_4
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_183_ net5 _076_ _042_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a21bo_1
X_252_ clknet_1_0__leaf_clk _026_ _010_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_235_ _073_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
X_166_ net2 VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__clkbuf_4
X_149_ _085_ _095_ _101_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__nand3_1
X_218_ _090_ _093_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__nand2_1
Xoutput17 net17 VGND VGND VPWR VPWR count[7] sky130_fd_sc_hd__clkbuf_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_251_ clknet_1_0__leaf_clk _025_ _009_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_2
X_182_ _040_ _041_ _110_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_234_ _073_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__inv_2
X_165_ _116_ _117_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__xnor2_1
X_217_ _068_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__clkbuf_1
X_148_ _096_ _097_ _100_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput18 net18 VGND VGND VPWR VPWR count[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_181_ _107_ _108_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_250_ clknet_1_1__leaf_clk _024_ _008_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_233_ _073_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__inv_2
X_164_ net10 _076_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__xor2_1
X_216_ net13 _067_ net2 VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_147_ _098_ _099_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__nor2_1
Xoutput19 net19 VGND VGND VPWR VPWR count[9] sky130_fd_sc_hd__clkbuf_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_180_ net19 net18 _076_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__o21a_1
X_232_ _073_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__inv_2
X_163_ _079_ _115_ _077_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_146_ net16 _074_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__nor2_1
X_215_ _086_ _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_129_ net7 _076_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_231_ _073_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__inv_2
X_162_ _081_ _084_ _113_ _114_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 ctrl VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_145_ net16 _074_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__and2_1
X_214_ _090_ _093_ _088_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ _080_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_230_ _073_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_161_ net8 net7 _076_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__o21ai_1
Xinput2 en VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
X_213_ _064_ _065_ net25 _032_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__a2bb2o_1
X_144_ net17 _074_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_127_ net8 _075_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_160_ _107_ _111_ _112_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__o21ba_1
Xinput3 rst VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_143_ net15 _074_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__xnor2_2
X_212_ _085_ _095_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__nor2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_126_ _077_ _078_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ _119_ _053_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nand2_1
X_142_ _087_ _090_ _093_ _094_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_125_ net9 _076_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_210_ _063_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__clkbuf_1
X_141_ net13 net12 _074_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_124_ net9 _076_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ net4 _091_ _092_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_123_ _075_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_199_ _053_ _096_ _054_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__o21ai_1
X_122_ _074_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_198_ net15 net14 _076_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_121_ net1 VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_197_ _085_ _095_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__nand2_1
X_249_ clknet_1_0__leaf_clk _023_ _007_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 net4 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_196_ _051_ _052_ net23 _032_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a2bb2o_1
X_248_ clknet_1_1__leaf_clk _022_ _006_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_2
X_179_ _039_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__clkbuf_1
Xhold2 net9 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_195_ _106_ _102_ _103_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__and3_1
X_247_ clknet_1_0__leaf_clk _021_ _005_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_4
X_178_ net7 _038_ _119_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3 net11 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_194_ _119_ _107_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__nand2_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_246_ clknet_1_0__leaf_clk _020_ _004_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_4
X_177_ _084_ _113_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__xor2_1
X_229_ _073_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 net18 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_193_ _050_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__clkbuf_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_245_ clknet_1_0__leaf_clk _019_ _003_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_4
X_176_ _037_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__clkbuf_1
X_159_ net6 net5 net19 net18 _075_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__o41a_1
X_228_ _073_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__inv_2
Xhold5 net12 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_192_ net19 _049_ _119_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__mux2_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_175_ net8 _036_ _119_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__mux2_1
X_244_ clknet_1_1__leaf_clk _018_ _002_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_158_ _108_ _109_ _110_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ _073_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
Xhold6 net14 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ _108_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__xnor2_1
X_174_ _080_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__xnor2_1
X_243_ clknet_1_1__leaf_clk _017_ _001_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
X_157_ net5 _075_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__xor2_1
X_226_ _073_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_209_ net15 _062_ net2 VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ _104_ _107_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__nand2_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_242_ clknet_1_1__leaf_clk _016_ _000_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfrtp_2
X_173_ _084_ _113_ _082_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_156_ net6 _075_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__xnor2_1
X_225_ net3 VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__buf_4
X_208_ _096_ _061_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_139_ net11 _074_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_241_ net3 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__inv_2
X_172_ _033_ _034_ net21 _032_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_224_ _119_ net20 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__xor2_1
X_155_ net19 _075_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_207_ net14 _076_ _053_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__a21boi_1
X_138_ net11 _074_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_171_ _079_ _115_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nor2_1
X_240_ net3 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_223_ _071_ _072_ net22 _032_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a2bb2o_1
X_154_ _102_ _103_ _106_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__a21o_1
X_206_ _060_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__clkbuf_1
X_137_ _088_ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_170_ _079_ _115_ _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_153_ _104_ _105_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__nand2_1
X_222_ _092_ _091_ net4 VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__a21oi_1
X_205_ net16 _059_ net2 VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__mux2_1
X_136_ net12 _074_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_152_ net18 _075_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__or2_1
X_221_ net4 _092_ _091_ _032_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__a31o_1
X_204_ _100_ _055_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__xor2_1
X_135_ net12 _074_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_151_ net18 _075_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__nand2_1
X_220_ _032_ net24 _069_ _070_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a22o_1
X_203_ _058_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__clkbuf_1
X_134_ _086_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput4 net4 VGND VGND VPWR VPWR count[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_150_ net17 net16 net15 net14 _075_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__o41ai_1
X_202_ net17 _057_ net2 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__mux2_1
X_133_ net13 net1 VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__xor2_2
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput5 net5 VGND VGND VPWR VPWR count[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_201_ _097_ _056_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__xnor2_1
X_132_ net14 _075_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput6 net6 VGND VGND VPWR VPWR count[11] sky130_fd_sc_hd__clkbuf_4
.ends

